���P      �!sklearn.neighbors._classification��KNeighborsClassifier���)��}�(�n_neighbors�K�radius�N�	algorithm��auto��	leaf_size�K�metric��	minkowski��metric_params�N�p�K�n_jobs�N�weights��uniform��feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�gender��SeniorCitizen��Partner��
Dependents��tenure��PhoneService��MultipleLines��InternetService��OnlineSecurity��OnlineBackup��DeviceProtection��TechSupport��StreamingTV��StreamingMovies��Contract��PaperlessBilling��PaymentMethod��MonthlyCharges��TotalCharges�et�b�n_features_in_�K�outputs_2d_���classes_�hhK ��h��R�(KK��h�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�_y�hhK ��h��R�(KM:��h�i4�����R�(KhCNNNJ����J����K t�b�B�L                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �t�b�effective_metric_params_�}��effective_metric_��	euclidean��_fit_method��brute��_fit_X�hhK ��h��R�(KM:K��h�f8�����R�(KhCNNNJ����J����K t�b�Bpj       �?                                      �?       @      �?                                               @              �?       @�&`��?���b��?      �?              �?        Zas �
�?      �?       @      �?       @       @                       @       @              �?       @�2���?�wX!�x�?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @nC��x�?����3w�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�፿Po�?@}m[&?                      �?      �?6��9�?              �?                                                                      �?      @�d�Q�ϰ?ƙ���?                      �?      �??���@��?      �?                       @                                                               @ e��h�?\Z ��n�?                                              �?              �?                                       @       @                       @ J�hY�?���f��?      �?                        v�'�K�?      �?       @               @       @       @       @                       @                ����`�?[�mG�Z�?                                ��V��?      �?       @      �?               @                       @       @              �?       @.�jL��?�9��gb�?              �?      �?        �z2~���?      �?              �?                       @                       @              �?       @J̖p���?v��`�?      �?      �?      �?        ���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?g�)L�ٲ?u�w@o�?                                ��Vؼ?      �?       @      �?                                                              �?       @F��s��?���pQ�?                                �V�H�?      �?       @      �?               @       @                       @      �?      �?       @Q�E�*�?��T+�5�?              �?      �?        �'�K=�?      �?       @      �?               @                                              �?      �?7w\I`��?D��'�?      �?                        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @1[�yj�?�Dv�8P�?                      �?      �?��ۥ���?      �?       @      �?       @               @       @               @       @               @
�R,�?���QQ^�?              �?      �?        6��9�?      �?       @      �?                                       @       @              �?       @3��l�?�e�˸�?      �?      �?      �?      �?�'�K=�?      �?              �?                                       @                      �?      �?*L����?kj����?      �?              �?        6���?      �?       @               @       @       @               @       @       @      �?       @J̖p���?R� (<��?      �?              �?              �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?E�(Ţe�?wk� ���?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?1[�yj�?���Lm�?                      �?      �?�6��?      �?                       @       @               @       @       @      �?              �?������?c�l^)s�?                                ��ۥ���?      �?              �?                       @       @               @              �?       @d�Q���?��=��?      �?                        ���V،?      �?              �?                                                              �?       @p�l�?=(����?      �?                        6��9�?      �?                                                               @              �?        ƽ�,u��?����<��?      �?                        3~�ԓ��?      �?       @      �?       @       @       @       @       @              �?              �?�Dz�rv�?�z*ՈD�?      �?              �?      �?�'�K=�?      �?              �?               @       @               @       @      �?      �?      �?�,���?�?�r �	��?      �?      �?      �?      �?��ۥ���?      �?       @      �?       @       @                       @       @              �?      �?����Z��?��-9y��?                      �?      �?{2~�ԓ�?      �?       @      �?                       @       @                              �?       @<��u�4�?z�;�9A�?      �?                        Zas �
�?      �?       @      �?       @               @               @       @              �?       @�(Ţe�?�4�1�?                      �?        ��V��?      �?                               @               @                      �?      �?      �?N��b��?�&�'�?      �?      �?                ?���@��?              �?                                                                      �?        ��Po��?nS�<�ǃ?              �?      �?        >�]���?      �?       @      �?       @       @       @       @                      �?               @�:��?���P�"�?              �?      �?                      �?       @      �?               @                       @                      �?       @���l	�?}����?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�0[�yjv?t������?      �?              �?      �?���@��?      �?       @                               @       @       @              �?      �?       @�7�B�]�?��D�5H�?      �?                                      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @���Z��?g�Ǘ��C?      �?      �?      �?        ���V،?      �?              �?                                                                       @cX�~k��?�#��Z�?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                       @#w\I`ޓ?��xIv?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                nC��x�?��ј��?      �?      �?                F���@��?      �?              �?                                       @       @              �?       @]�F�?+ߙ�v�?      �?      �?      �?        ��RO�o�?      �?       @      �?               @       @                       @              �?       @X~PT��?�I�Bf�?                      �?      �?�ԓ�ۥ�?      �?       @               @                       @                       @              �?�o��z�?�;-�	��?                      �?        SO�o�z�?      �?       @      �?                       @       @                              �?      �?>�� Q��?g!ի�g�?                                              �?       @      �?                                                              �?       @��8j��?g1'+<�z?      �?                        Zas �
�?      �?              �?                                                              �?      �?��j1v�?g��*��?              �?                              �?              �?               @                                              �?       @�HT�n�?�4]0#�y?                      �?      �?$Zas �?      �?               @      �?      �?      �?      �?      �?      �?                       @��N�ԑ?�g�x���?                                6��9�?      �?              �?               @       @                              �?               @���w��?��Yc(�?                                �@�6�?      �?              �?                                       @       @              �?       @� 6\.2�?����ɩ?      �?                                      �?              �?                                                              �?       @X-�r�?�3�
'x?                                3~�ԓ��?      �?       @      �?                       @               @       @              �?       @�^<��u�?g��q}�?      �?              �?      �?�K=��?      �?              �?               @       @       @       @       @       @                3��g�?�q���d�?      �?                        ���@��?      �?       @      �?       @       @       @       @       @       @      �?              �?�L�cX��?�=G�P�?      �?              �?        6��9�?      �?       @      �?                                               @              �?       @UUUUUU�?�D����?      �?                        {2~�ԓ�?      �?                                               @                              �?       @��x�]��?PD*����?      �?              �?        �@�6�?      �?              �?               @       @                       @              �?       @�jL�*�?�8�|�B�?      �?              �?      �?!�
���?      �?                       @                       @       @       @      �?      �?        m$���?L���+'�?      �?              �?      �?SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����`�?�?�)�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @,1[�yj�?`Ĭ)�?              �?                �]�����?      �?       @      �?                                                              �?        �u�b���?������?              �?                �'�K=�?      �?       @      �?                       @               @       @                       @�^<��u�?R�#M��?                      �?      �?�ԓ�ۥ�?              �?               @               @                       @       @      �?      �?�7�B�]�?go��׸�?      �?                                      �?                                                                              �?      @2NaJ̖�?�i)��h?      �?                        �K=��?              �?                                                                      �?        ?�]�FR�?�� O��?                      �?        �
��V�?      �?              �?       @                               @       @      �?      �?       @&���[�?莂w�i�?              �?      �?        ���@��?      �?       @      �?               @                       @                      �?       @��r�9�?X�i��?      �?              �?      �?�'�K=�?              �?               @                                                      �?        FaJ̖p�?ޚL�
��?      �?              �?      �?�@�6�?      �?       @               @                               @                      �?        �������?n��д?                                $Zas �?              �?                               @               @       @              �?      �?�{B���?`�Fb���?                      �?      �?>�]���?      �?       @               @       @                               @      �?                ����`�?B�9��	�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?        �U�����?qpTV�?      �?              �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @               @���T��?L��'���?      �?                         �
���?      �?              �?               @                       @                      �?       @�@��~�?K`K�Im�?              �?      �?        ���Vج?      �?       @      �?                                                              �?       @,�����?�J�Tt��?      �?              �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����`�?c%��ި?      �?                              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ��w����?3��)f��?                                P�o�z2�?      �?       @      �?       @       @               @       @       @       @              �?mZq�$K�?���Wl��?                      �?      �?!�
���?              �?               @                       @                       @                ��"X~P�?�ųR	�?      �?              �?        �z2~���?      �?              �?               @                               @              �?      �?H*��E�?�QI���?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @��N�ԑ?�Ր�,u?      �?                        �ԓ�ۥ�?              �?                               @               @       @                       @��̱���?nB�C7��?      �?      �?      �?        6��9�?      �?                       @               @               @                                �w�ӥ��?�)M���?                                �K=��?      �?              �?                                                              �?      �?�¯�Dz�?��z"Z��?                      �?        �'�K=�?      �?                       @                       @               @       @              @��@���?d�?���?      �?              �?        �6��?      �?       @                               @       @               @      �?              �?�돗�(�?'��]V��?      �?              �?        �6��?      �?               @      �?      �?      �?      �?      �?      �?       @                ���C�?���}h�?                                Zas �
�?      �?       @               @               @       @       @       @       @              �?�WH�%��?�vu
�?      �?              �?      �?              �?              �?                                       @       @                      @��Y;��?PK�h"��?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @����[�?+T�ʟ?      �?              �?      �?ܥ���.�?      �?                               @       @                              �?      �?      �?ͤ=����?�1s�p�?      �?              �?        {2~�ԓ�?      �?       @                       @               @       @              �?              �?L�*g��?�̖fVp�?      �?              �?      �?[as �
�?      �?       @      �?       @               @       @                                       @}�mu��?�cFۣ��?                                �ԓ�ۥ�?      �?       @      �?                                       @                      �?       @�WH�%��?["$NK;�?      �?              �?      �?�ԓ�ۥ�?      �?       @               @       @       @       @                       @      �?      �?�Kn��4�?�'.�Y@�?                              �?�K=��?      �?       @      �?               @               @       @       @       @      �?       @'Y��M�?KPULD��?              �?                �]�����?      �?                       @               @       @               @              �?      @����e�?���f��?      �?                        �]�����?      �?       @      �?                                               @                       @�{B���?��7�sL�?      �?                        ��RO�o�?      �?       @      �?                                       @                                b�(Ţe�?~S��f��?                                F���@��?              �?                       @                                              �?       @|+�oM�?���E�g�?                      �?      �?�]�����?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��N�Ա?���b���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      �?�፿Po�?fN
u�w*?      �?              �?      �?      �?      �?       @      �?               @       @               @       @       @      �?       @�p���?��o��'�?      �?                              �?      �?       @                       @       @       @       @       @       @      �?        ffffff�?�G����?      �?              �?        �RO�o��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �^W-��?L�e��?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?                -h#���?=w���?                              �?��Vؼ?      �?                                       @       @       @       @              �?      @�%��f�?T�����?                      �?        ��RO�o�?      �?              �?                               @       @       @      �?      �?       @U:'>���?�W����?      �?                        �D+l$�?              �?                                       @       @       @              �?       @Ͽk�.M�?�y6>�?      �?              �?        �ԓ�ۥ�?      �?       @                       @               @       @              �?      �?       @�돗�(�?�V�j���?                                F���@��?      �?              �?               @                                      �?      �?      @�k�.M��?����?                      �?        �z2~���?      �?                                       @       @                                       @���@���?�0�����?                                3~�ԓ��?      �?       @      �?       @       @       @               @       @                      �?�1���?F���z��?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�%��}�?D�28�I�?      �?              �?      �?�'�K=�?      �?       @               @                       @       @              �?                b����,�? $NK;��?      �?              �?      �?�]�����?      �?       @                               @       @       @       @      �?      �?      @���Y;�?AW(j�K�?                      �?      �?      �?      �?       @               @       @       @       @               @       @                B�/����?M�(�bp�?      �?              �?      �?��ۥ���?      �?              �?       @       @       @       @       @               @              �?:'>���?sS���?      �?              �?        F���@��?              �?               @       @                                                      @��"X~P�?-V�a�?      �?      �?      �?        e�v�'��?              �?                                                                      �?        �?���,S��?              �?                ��RO�o�?      �?              �?       @       @               @               @      �?      �?      @��C���?�K ��'�?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?D�2� Ѝ?                                                      �?                                                                               @_����,�?W�n�X�E?              �?      �?        ���V،?      �?              �?                                                              �?       @1�L�5A�?8v\l�?      �?                        �@�6�?      �?                       @                                       @              �?        ��_���?�"�1Ȣ?                      �?        ���V،?              �?                                               @       @                       @X�ڙ���?������?                                3~�ԓ��?      �?       @               @       @       @       @       @               @      �?      �?��*��?������?              �?                H���@��?      �?       @      �?               @                               @              �?       @+�oM��?�aW�@�?                                �
��V�?      �?                       @                       @                      �?              @����?+P�͏�?      �?              �?        �D+l$�?              �?                                               @       @              �?       @2NaJ̖�?[��;��?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                      @1[�yj�?�4b�9��?                                ?���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�k�.M��?�B�2�?                      �?                      �?               @      �?      �?      �?      �?      �?      �?              �?        �'�F7�?O���&?      �?                        3~�ԓ��?      �?              �?       @       @       @                       @              �?      �?�o2���?bJ�U$��?                                (�K=�?      �?                       @               @       @       @       @       @                4�G�Ɉ�?��q���?      �?                        �'�K=�?      �?              �?                                                                        ���S��?���u���?      �?              �?      �? �
���?      �?                                       @                              �?              @���7q�?fO�M̶�?              �?                $Zas �?      �?              �?                                               @              �?       @h#���?��g$�i�?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?�d�Q�ϐ?'�d��+\?      �?              �?      �?$Zas �?      �?                                       @                                      �?       @�7q���?�����4�?      �?              �?      �?SO�o�z�?              �?                       @       @                       @      �?      �?      �?����7�?�v�A���?      �?              �?      �?ܥ���.�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �%��f��?5����?                      �?      �?�RO�o��?      �?       @      �?       @       @                       @              �?                Q�E�*�?i�$d�?                      �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �L�5A �?�ϖ��?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?       @       @                                              �?      �? ʣ��8�?�tdlK�?      �?                        ��V��?      �?       @      �?               @       @               @       @       @              �?����Z��?�S��Vk�?      �?              �?        6��9�?      �?       @      �?       @       @               @                              �?      �?r�9ֳv�?�0�"ml�?      �?      �?      �?        �z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�bѲ
n�?1Q��a�?      �?                        ,l$Za�?      �?                       @                       @       @              �?               @}�mu��?+��G
Z�?      �?                        ���V،?              �?                                                                              @�c=kgҮ?��0A�b?              �?                �ԓ�ۥ�?      �?       @      �?       @               @       @       @       @       @              �?mZq�$K�?�N+OT��?                                �6��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @n��W�?N�9�z�?      �?                        >�]���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�j1v�?10qum�?      �?                        6��9�?      �?                                                                              �?       @O�0@�b�?"u�m묦?              �?      �?        (�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?      �?X��M+�?(�5�l�?                                �ԓ�ۥ�?      �?                       @               @       @       @       @       @      �?      �?���7q�?g\�8�q�?      �?              �?      �?Zas �
�?      �?                       @       @                                      �?      �?      @V:'>���?q�s��ȸ?              �?                F���@��?      �?       @      �?                                               @              �?       @��-�jL�?Y���_�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @9�%��}�?V���+�?                              �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�k�.M��?CB+��?      �?      �?      �?        �z2~���?      �?              �?                                       @       @              �?       @��ǰ2��?uk:���?      �?              �?      �?�ԓ�ۥ�?      �?       @                       @       @       @       @       @       @      �?        9�WH�?� �P@��?      �?              �?        �K=��?              �?               @       @               @               @       @      �?        �������?�txn���?      �?                        �ԓ�ۥ�?      �?       @      �?                                                                      @!�����?z~0�t5�?              �?      �?        $Zas �?      �?              �?                                       @       @      �?      �?        �jL�*�?_���0�?      �?              �?      �?$Zas �?              �?               @               @       @                       @      �?      �?�!�����?V�0��ӷ?      �?              �?      �?      �?      �?       @      �?                       @                       @       @      �?      �?�?y4��?�����?                                p�z2~��?      �?       @      �?       @               @               @              �?              �?p2��g�?���J
��?      �?                        SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?      �?                -h#���?�0dA"��?                      �?      �?�
��V�?      �?              �?                                               @              �?       @O�)���?��O�?      �?                        �D+l$�?      �?              �?       @       @       @                                      �?      �?�H*���?D�����?                                              �?               @      �?      �?      �?      �?      �?      �?                      @���C�?ݘ<$3(?      �?                        �ԓ�ۥ�?      �?              �?                               @                              �?        �8�)1[�?F��� �?                      �?        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @E�(Ţe�?4}����?                                �]�����?      �?               @      �?      �?      �?      �?      �?      �?              �?      @n��W�?�7�!\��?      �?                        ���V،?      �?              �?                                                                      �?���S��?�s�1�Ό?      �?                        ?���@��?      �?                               @               @       @                      �?        -�Q����?7,{Hʁ�?                      �?        (�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?m+�oM�?�4�O�W�?      �?              �?      �?      �?      �?       @               @       @       @       @       @               @      �?        B�/����?Ÿ h�?      �?      �?      �?        6��9�?      �?       @      �?                                               @              �?       @��ds��?��|!.��?      �?              �?      �?�ԓ�ۥ�?      �?       @               @               @       @       @       @       @                }x�/���?�a$Y���?      �?                      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?                      �?�r@��?���@7<�?      �?                      �?[as �
�?      �?       @                       @               @       @       @      �?      �?      @�ti��|�?������?                                ?���@��?      �?              �?                                                                       @�V�ߚ�?��oy��?      �?                                      �?                                                       @                      �?      @��Dz�r�?�	�fp?      �?              �?        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?                -h#���?uD{@O��?      �?                              �?      �?       @      �?               @       @               @       @      �?      �?       @�e� ��?��ҡ���?      �?      �?                �]�����?      �?       @      �?                               @       @                      �?        ]�F�?�P��L��?                                $Zas �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @nC��x�?��=��?      �?                        !�
���?      �?       @      �?               @       @       @                              �?       @X�~k� �?'��r�?                                �ԓ�ۥ�?      �?       @      �?                               @       @                      �?       @�p��R�?��V
u��?      �?      �?      �?      �?v�'�K�?      �?       @      �?               @       @       @       @       @      �?      �?       @��l��?�W�φ�?      �?              �?      �?SO�o�z�?      �?       @               @       @                       @                      �?        �A6w\I�?�p�r�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @��N�ԑ?n�CT�?      �?                        �6��?      �?       @      �?                       @       @       @              �?                ���`p�?��:}�?                                              �?              �?                                                              �?       @�c9�?o��W�w?      �?              �?        ��RO�o�?              �?                       @       @       @       @       @      �?      �?       @��V���?�Ni0�`�?                      �?        3~�ԓ��?      �?              �?       @               @                              �?      �?      �?�b��!�?���b�8�?      �?              �?      �?F���@��?      �?                       @                                              �?      �?       @[�՘H�?L6�u�v�?                              �?�'�K=�?      �?              �?                                                                        �돗�(�?&C���Լ?      �?                        !�
���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @��w����?,j&-3��?              �?      �?        F���@��?              �?                                               @       @                       @�����9�?��a�?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?                      @F��1��?��ֺ�?                                �o�z2~�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?����[�?�����Q�?                      �?        �ԓ�ۥ�?      �?                               @               @                                       @��f��?���d!6�?                                              �?              �?               @                       @                               @�H*���?���l�~?                      �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @8�]�FR�?�R�ʵ?      �?              �?      �?F���@��?      �?                                                                                        q%�yO��?�Ea�x�?                      �?        �@�6�?      �?              �?                       @       @                      �?               @��.h�?��I}u�?      �?                      �?��.�d��?      �?       @               @       @               @       @       @       @      �?      @Ͽk�.M�?=���h�?      �?              �?      �?�]�����?      �?                       @               @       @       @       @       @      �?      �?Y���d�?P��~3�?      �?                        ���V،?              �?                       @       @       @                              �?      �?�~k� 6�?2_�\H�{?      �?                        Zas �
�?      �?       @      �?               @                                              �?      @��r�9��?�e�qE+�?      �?              �?        >�]���?      �?       @      �?               @                       @       @      �?              �?��'t �?��b���?      �?              �?      �?�RO�o��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�፿Po�?#��w��?      �?      �?      �?        p�z2~��?      �?       @      �?       @                                                      �?       @���Z�K�?�w�i+��?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�L�5A �?4Uo����?      �?              �?        �z2~���?      �?                       @                                       @              �?        V�&#��?��I�L}�?      �?                        �o�z2~�?      �?       @      �?       @       @               @               @      �?               @�������?r:��Y
�?                      �?      �?�D+l$�?      �?       @               @       @               @                      �?              @��@���?r�|�8��?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                      @]����`�?)�Fw�?      �?              �?      �?��V��?      �?       @      �?       @       @       @       @                       @              �?�0%fK�?��}`�?      �?                        ���V،?      �?              �?                                                                      @���S��?d��"�?      �?              �?        H���@��?      �?       @      �?       @       @                       @                      �?        m��W�?f�R�qh�?      �?      �?      �?        �6��?      �?       @      �?               @       @               @       @              �?       @�+$����?�m.Gx�?      �?                                              �?               @                                                              @P��*�?��a���T?                      �?        ��ۥ���?      �?       @      �?       @       @                       @              �?              @�:��?�y�� @�?                              �??���@��?      �?       @      �?               @                       @                              @�=����?e4jd~�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?�t&���P?      �?              �?      �?��ۥ���?      �?       @      �?       @       @       @       @       @       @       @      �?        �:]��#�?b�8K��?      �?                        �D+l$�?      �?       @      �?                               @               @              �?      �?8�B�]��?�S�����?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @Y�)L�ْ?CX�?|Ͳ?      �?              �?        �RO�o��?      �?       @      �?               @       @               @                      �?       @d�#�6��?�TQ�#�?                              �?�K=��?      �?       @      �?       @       @       @       @       @       @       @      �?      �?]�FR,�?`{�D~�?                      �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?                1[�yj�?_�VP��?      �?                      �?	��V��?      �?                               @       @       @       @       @      �?               @B�/����?%�y\�?      �?                        ��Vؼ?              �?               @               @       @               @      �?              @]<��u��?���,�G�?                      �?      �? �
���?      �?              �?       @       @                                                       @9�WH�?ƕ]7L�?      �?      �?                ��.�d��?      �?       @      �?                                                              �?        �}��j�?Ak�5%�?      �?              �?        !�
���?      �?       @      �?       @               @       @       @       @      �?      �?       @@�MF��?�b
��?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�%��}�?����?      �?              �?      �?              �?              �?                                       @       @              �?       @C)-���?X�dޛـ?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�፿Po�?��Š���?      �?              �?        �D+l$�?      �?       @      �?       @       @       @               @       @      �?      �?       @�ć7�B�?6�����?      �?      �?                �@�6�?      �?       @      �?               @       @               @       @              �?       @}䛌8j�?�̡��?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @���C�?d1G���?                                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @$�$0�	�?���ݕU�?                                              �?       @      �?                                               @              �?      @b�(Ţe�?;�
���?                                ܥ���.�?              �?               @       @                       @                      �?       @q%�yO��?�Hվ���?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @-h#���?���M�r?                                ?���@��?      �?       @      �?               @                                                        ���J�?"�Wi�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @E�(Ţe�?���ܧ?      �?              �?      �?�K=��?      �?       @               @               @               @       @       @      �?       @�j1v��?��z�?                      �?        Zas �
�?      �?       @      �?               @                       @       @       @      �?        /��:]�?f�)���?      �?                        ���.�d�?      �?       @                       @       @       @       @       @       @              �?&�1�L��?�hP����?      �?              �?      �?��Vؼ?      �?              �?               @               @       @       @              �?       @���?$�jg�;�?              �?      �?        ��V��?      �?       @      �?       @               @               @       @                        5&����?2v͔o��?      �?              �?        6��9�?      �?       @               @               @               @       @      �?              @�I�:Bl�?�؋��]�?                      �?      �?�ԓ�ۥ�?              �?                                       @       @              �?              @-����?AF͙(�?      �?      �?                              �?       @      �?                       @               @                      �?       @r�9ֳv�?.v&����?      �?              �?        ��RO�o�?      �?                               @       @       @       @       @       @              @9�WH�?P�?�\-�?      �?              �?      �?      �?              �?               @       @       @       @       @       @       @      �?      �?1�z�Τ�?E~�[�?              �?                ���V،?      �?       @      �?                       @                                      �?       @333333�?��L�?              �?                ���Vج?      �?              �?               @                       @                      �?       @��a�(�?F͙(�?      �?                        �]�����?      �?       @      �?       @                               @       @              �?       @��¯�D�?9� o���?      �?              �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?-h#���?���L�z�?      �?              �?      �?p�z2~��?      �?       @      �?               @                       @       @              �?       @E������?�pȝw�?                      �?        H���@��?      �?              �?                       @                                      �?       @����9��?-{-�F�?      �?                                      �?                       @                                                      �?      @ئ�N��?X2��3n?      �?              �?      �?!�
���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�?"K�}���?                              �? �
���?      �?       @                                                                      �?      @�F���?o�+J�j�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?�^/��"?      �?                        e�v�'��?      �?       @      �?               @                                              �?        ��*��?��B ���?                      �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @E�(Ţe�?=���o�?                      �?      �?Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @ò
n�ͭ?e>�?أ�?      �?                      �?���V؜?      �?       @      �?                       @                       @                       @�፿Po�?0��g�&�?              �?                ���Vج?      �?              �?                                                              �?      @b����,�?QSU봡?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @����'t�?��ʲ?                                �@�6�?      �?                       @       @                                                      @�a/��?�7��w��?                                ��RO�o�?      �?              �?               @       @       @               @      �?      �?      �?�Gm?C�?�5-N(��?      �?                              �?      �?       @               @       @       @       @       @       @       @                :Blӊ{�?� Ȣ0l�?                      �?      �?��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @Xph>ׯ?WSѭJP�?      �?      �?      �?        ��V��?      �?       @      �?                                       @       @              �?       @V�;�RG�?������?      �?                        �ԓ�ۥ�?      �?       @               @       @       @       @               @      �?      �?      �?��'�F7�?��<����?      �?                                              �?                                               @       @              �?      @�����9�?���W�i?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?               @       @               @       @       @      �?       @e0
84��?8�����?      �?                        ��Vؼ?      �?                                                                              �?      @?y4���?��	_u�?                                ?���@��?      �?              �?                                               @              �?       @Y���d�?�I$a��?                                (�K=�?              �?               @               @       @       @       @       @      �?        �n�)L��?7GUo���?                              �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @F��1��?Y��N��?      �?              �?      �?�z2~���?      �?                       @                       @                      �?              �?~�ɣ���?��o��?                      �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?-h#���?�{NN�c�?      �?              �?        ��RO�o�?      �?                       @                                              �?              �?Y���d�?���ڸ�?      �?                        �K=��?      �?               @      �?      �?      �?      �?      �?      �?                      @^��Z��?al� g�?      �?      �?      �?        �K=��?      �?                       @       @               @                      �?      �?        ��8�)1�?úy�H�?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?                       @]����`�?���0��?                                �@�6�?      �?                                                               @              �?       @jL�*g�?9�S' �?                      �?      �?Zas �
�?      �?              �?               @       @               @                      �?      �?[ݧ����?Z~�����?      �?                      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @#w\I`ޓ?,�q��̂?              �?      �?        ��ۥ���?      �?       @               @       @       @       @               @       @      �?        v�z��?��b{v�?                                v�'�K�?      �?       @      �?       @       @       @       @               @              �?        o��T�?��9�H�?              �?      �?        �
��V�?      �?              �?                       @       @       @               @              �?r�9ֳv�?v�����?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        	�Y e�?U`(G:<�?      �?                        �V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @                n��W�?;d��"�?                      �?        ���.�d�?      �?              �?       @               @               @       @       @      �?        �$K!��?b�0TKy�?                      �?        ��RO�o�?      �?              �?       @       @               @       @       @      �?              @�<5���?i�m�d��?      �?      �?                �@�6�?      �?       @      �?               @       @       @       @       @              �?       @��o2��?�w�@G2�?      �?      �?      �?        �]�����?      �?       @      �?               @                       @       @              �?       @mӊ{'Y�?����"�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?      @1[�yj�?G���>[f?      �?              �?      �?�'�K=�?      �?                                       @                                      �?       @�'�F7��?%<^9i�?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�፿Po�?QSU봑?      �?                        ��Vؼ?      �?                       @               @       @               @              �?        _ph>��?7WK�|�?      �?                      �?$Zas �?              �?               @                       @       @              �?                �?j�-�+�?                              �?�z2~���?      �?                                               @                      �?      �?       @5w\I`��?���=jA�?                      �?                      �?              �?                                                              �?      @�A6w\I�?����w?      �?      �?      �?        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?0�'Tn'�?      �?                        �@�6�?      �?       @      �?                                                              �?       @E_r[ݧ�?������?                                ��V��?      �?       @      �?               @               @       @       @      �?      �?        )���G��?���`���?      �?                        �K=��?      �?                                               @                       @                �Po���?�L/=��?      �?              �?        >�]���?      �?              �?                                       @       @                      @+�oM��?Ⱥ��D8�?              �?                ?���@��?      �?       @      �?                                       @       @              �?       @J�hY7�?l)-�e��?      �?      �?      �?        ,l$Za�?              �?                       @                                              �?       @�c=kgҾ?�oN�:��?      �?              �?              �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?^��Z��?;e��k��?                      �?        p�z2~��?      �?       @      �?                       @               @       @              �?       @����e0�?�����O�?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?��f��}�?M'�1m�?      �?                                      �?                       @                       @                              �?       @g{����?��4�p?      �?              �?        >�]���?      �?              �?                                               @      �?      �?       @m$���?[���r��?      �?              �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                       @����[�?;����?      �?              �?        SO�o�z�?      �?       @      �?                       @       @       @       @              �?        �g{���?7�m��?      �?                      �?��ۥ���?      �?       @      �?       @       @                                      �?      �?      �?b�(Ţe�?H�mj1�?                                �V�H�?      �?              �?               @       @       @       @       @       @      �?        A���Kn�?�o�/
�?      �?                        ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?m+�oM�?������?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @�Y;���?ZX�ħJr?                      �?        �
��V�?      �?               @      �?      �?      �?      �?      �?      �?                      @���@��?�Ǘ���?      �?              �?              �?              �?               @       @       @       @       @       @       @      �?       @&��f���?�A��t�?              �?                �@�6�?      �?              �?                       @       @       @       @      �?      �?        �ht3Na�?��'&���?              �?      �?        p�z2~��?      �?       @      �?                                       @       @              �?       @������?(Z���?      �?      �?      �?        F���@��?      �?              �?               @       @               @       @              �?       @�M+�d�?�.x%}�?                      �?      �?�
��V�?      �?       @      �?       @                               @       @      �?              @�=�� Q�?�.���?      �?              �?        �D+l$�?      �?       @                                                                               @���'�??��<�?                      �?        �V�H�?      �?       @               @                                                                jL�*g�?�΅D�!�?      �?      �?                �z2~���?      �?       @      �?               @       @               @       @              �?       @�]�FR�?)pl�3�?                                F���@��?      �?              �?                       @               @       @              �?       @KS}䛌�?e�����?      �?      �?                �K=��?      �?       @      �?                       @               @       @              �?      �?�)1[�y�?.�P�1�?                      �?      �?6��9�?      �?                                       @       @                                      �?��J�ć�?\����?                                 �
���?      �?       @      �?                       @                                      �?       @�AQ�s��?{��Î�?      �?      �?      �?        F���@��?      �?       @      �?                                                              �?       @/M��o2�?9���a�?                                F���@��?      �?                                               @       @       @              �?      �?L�*g��?O�I���?                                P�o�z2�?              �?                       @               @               @                       @�=�� �?竬���?                      �?        �'�K=�?      �?              �?                                       @       @                       @�E�*�A�?�P{�C�?                      �?      �??���@��?      �?       @                       @               @                              �?      @/�Q���?浚��X�?      �?                        �z2~���?      �?       @      �?                               @       @                      �?       @���l	�?�MXo�l�?      �?              �?      �?H���@��?      �?              �?                                       @       @      �?      �?       @���T��?~�;v���?      �?                        ��Vؼ?      �?       @      �?                                                              �?       @
n��W�?�>c��ٴ?              �?                $Zas �?      �?       @                                                       @              �?      @�e� ��?1Q��a�?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?       @#w\I`ޓ?6��pq?              �?      �?        	��V��?      �?       @      �?                                       @       @              �?       @����_��?h�wp��?      �?                        ��V��?      �?              �?               @               @                       @                r�g�L��?3��p�?                      �?        6��9�?      �?       @      �?       @               @       @               @      �?      �?       @�O�n��?(z����?      �?                                      �?                                                                              �?       @ꏗ�(��?��ׇh?                              �?6��9�?      �?       @               @       @               @       @                      �?      @�8�)1[�?p:��Y
�?              �?                $Zas �?      �?       @      �?                       @               @       @              �?       @^��C��?�c�A��?      �?              �?        p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?                       @���6�?�g�x��?                                �@�6�?      �?                                               @                              �?        ]<��u��?wm��П?      �?              �?      �?Zas �
�?      �?       @      �?       @       @                       @       @      �?      �?       @�*g���?�n���?                                �'�K=�?              �?                       @                                              �?       @}�mu�?��V齸?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                      @��N�ԑ?'u��&[�?                      �?        	��V��?      �?       @      �?                                       @       @                       @_��"s��?��c��?      �?              �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����'t�?��8��?      �?              �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @���6�?�-1��?      �?                        �6��?      �?       @      �?       @       @                       @       @      �?      �?       @�+$���?�չ��?      �?                        v�'�K�?      �?       @      �?               @                               @                      �?��%���?H+s6 �?                      �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�፿Po�?#���뤛?      �?              �?      �?���V،?      �?              �?                                       @       @              �?        �r�9ֳ�?]�i�#��?                      �?      �?�ԓ�ۥ�?      �?                       @                       @                      �?      �?        䶺O_�?֋��?                      �?        >�]���?      �?              �?       @       @       @               @       @      �?      �?      �?������?)ܼ�V�?              �?      �?        �'�K=�?      �?       @      �?                       @       @                              �?       @�{B���?Ȧ���N�?                      �?        P�o�z2�?              �?               @               @               @       @      �?      �?       @ J�hY�?��Lj\�?              �?      �?        ��ۥ���?      �?       @      �?       @       @       @       @                       @      �?      �?�*���?�����?      �?                        �@�6�?      �?                       @               @               @                                �3��x��?�� ����?      �?              �?      �?�K=��?      �?       @      �?       @       @       @               @       @      �?      �?       @o��z���?~=,`��?              �?      �?        ���@��?      �?       @      �?               @       @               @                      �?       @����'t�?s�����?              �?                ���V؜?              �?                                                                               @�k�.M��?p&���{?                      �?      �??���@��?      �?                               @               @                                      @&���[�?/�9��?      �?                        �'�K=�?      �?       @      �?                                       @       @              �?       @Τ=����?��%�q�?      �?              �?              �?      �?       @      �?               @       @       @       @       @       @      �?       @-�<5��?�]����?      �?                        �V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @               @8�]�FR�?����S=�?              �?                �'�K=�?      �?       @      �?                                                              �?       @�ئ�N�?�z�Z�Z�?                                3~�ԓ��?      �?       @      �?               @       @               @       @      �?      �?      �?�#�d�Q�?����`�?      �?      �?                p�z2~��?      �?       @      �?               @                       @       @              �?       @;�RG�m�?�C9���?      �?                        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @                8�]�FR�?UO���?                                ���V؜?      �?              �?               @                       @       @                       @r@���?���5�?                      �?      �?��ۥ���?      �?                       @       @       @       @                       @              �?S��*�?M��a��?      �?              �?        �K=��?      �?                       @       @               @               @       @      �?      �?�c9�?NY:�Z.�?      �?              �?      �?�@�6�?      �?              �?                                       @       @                       @���l	�?��C���?              �?                ���V؜?      �?              �?                       @               @                      �?       @�������?'��?      �?                        �'�K=�?      �?              �?                                                              �?      @cX�~k��?��b�v�?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        E�Ή�?|yw�;�?      �?                        ���V،?      �?                       @                                                      �?       @�0@�b��?��UR�g�?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?�o��'�r?                                v�'�K�?      �?                       @       @       @                               @      �?        �#�d�Q�?���$���?      �?              �?      �?��RO�o�?      �?                       @       @                               @       @      �?        �o��z�?��%J]��?                                �z2~���?              �?                       @       @       @       @       @      �?               @�L�5A �?4\���f�?      �?              �?        ?���@��?              �?                       @                       @       @              �?       @���Z�K�?�5X��?              �?                      �?      �?       @      �?       @       @       @       @               @       @      �?        �4�u�b�?��n&��?      �?      �?                ��ۥ���?              �?               @       @                       @       @      �?      �?       @�<݌S�?�D5�/K�?                      �?        ��V��?      �?                       @       @       @                       @       @                ������?��y�� �?      �?                        H���@��?      �?              �?                                                                       @����e�?����C�?                      �?        !�
���?      �?                       @       @               @                      �?      �?        ����?D�6���?              �?      �?        v�'�K�?      �?       @                       @       @               @              �?      �?        �9�፿�?���4�m�?                      �?      �?��V��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�^W-��?�:�	�?      �?                        p�z2~��?      �?                                       @                                      �?      @�b��!�?��d���?      �?      �?                e�v�'��?      �?                                       @       @               @      �?                ��M+��?�ڸd4��?      �?              �?      �?F���@��?      �?                                                       @       @      �?      �?       @�1����?5��\�?                      �?      �?6���?      �?              �?               @       @               @                      �?       @^!ї�V�?|��iH�?                      �?        H���@��?      �?       @               @       @       @                       @      �?               @NF���?I։���?                      �?         �
���?      �?       @               @       @       @       @       @       @      �?      �?      �?C)-���?�=�i���?                      �?        �z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�6��w�?��G�?                      �?        ��V��?      �?       @      �?       @       @               @       @              �?      �?        w\I`��?�nZv�?                      �?        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @�X����?/�,H��?      �?                        ���V؜?              �?                                                                               @��w����?J-�v?      �?                        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�d�Q�ϐ?.W�ж?              �?                ,l$Za�?      �?              �?               @       @                       @      �?              �?��Y;��?(bmweU�?                      �?        ��Vؼ?      �?              �?                       @                                      �?        �ئ�N�?��U�Ҳ?      �?              �?      �?��ۥ���?      �?                       @       @                                      �?              @B����? ���^�?      �?              �?        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @,1[�yj�?��(�X�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?��J�iҡ?              �?                ��V��?              �?                       @       @               @       @       @      �?        ��Dz�r�?���?l��?                      �?        ��ۥ���?      �?       @               @       @       @       @       @       @       @               @C)-���?�&���;�?      �?              �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @              �?8�B�]��?�T�1��?      �?              �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @      �?      @�`ph>�?�yofC�?                      �?      �?                      �?               @                                                                �e0
84�?Vp���V?                                �z2~���?      �?                                                                              �?       @�?=o�v˭?                      �?        ���V،?      �?                                                                              �?      �?X�ڙ���?@f3­/}?                                ?���@��?      �?              �?                                       @                      �?       @T�n�W�?.�:��̠?                      �?      �?�z2~���?      �?       @      �?       @       @                       @       @              �?       @���Kn��?/�8S]f�?                      �?              �?      �?       @      �?       @       @       @               @               @                H���<�?9�
�!�?      �?                        �K=��?      �?       @      �?       @       @       @       @       @       @      �?              �?�e0
84�?�����?      �?              �?        SO�o�z�?      �?       @      �?       @               @                       @              �?       @�FR,?�?+:��|��?                                �'�K=�?              �?                                       @                              �?       @���"X~�?�ގ�%κ?      �?      �?      �?        ���V؜?      �?       @      �?                                       @       @              �?       @�q%�yO�?	>��Ϟ?      �?                        [as �
�?      �?              �?                       @       @       @       @       @                �E�X���?<��!��?      �?                                      �?                                                               @              �?       @
84���?��nh:q?              �?      �?        �o�z2~�?      �?       @      �?               @       @               @              �?      �?      �?�6��`�?/ٴ���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @��N�ԑ?�rm[&"?                                	��V��?      �?       @                               @       @       @                      �?      @�돗�(�?c≋�?      �?                        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        n��W�?��g���?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�'�F7�?O���&?      �?              �?      �?�
��V�?      �?       @      �?       @       @                       @       @      �?               @)����?_X���?                                              �?       @      �?               @                                              �?      @Y���d�?����G�|?                      �?      �?ܥ���.�?      �?              �?       @               @               @       @      �?      �?        �;�$0��?��M[1O�?              �?      �?        �ԓ�ۥ�?      �?       @      �?               @               @       @       @       @              �?��Ͽ�?I.�0\��?              �?                SO�o�z�?      �?       @                               @                                               @;�^!��?l[g���?                                                      �?                                                                      �?      @\��r�?H��W�G?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @Y�)L�ْ?�Ǘ��c?              �?      �?         �
���?      �?              �?               @                               @                       @Ô�-�<�?�BY�3��?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�d�Q�ϐ?��3��c�?                      �?      �?�]�����?      �?       @      �?                       @                       @              �?        ����_��?��i>���?      �?                                      �?              �?                                       @                      �?       @q
Sb���?C7���|?              �?                              �?              �?               @                               @              �?       @�6��w��?�?Y�?                      �?      �??���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?�l��{3{?      �?                                      �?                               @                                              �?      @��"X~P�?�Ŏ���m?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @����[�?/(;p&k$?                      �?      �?      �?              �?               @       @       @       @       @       @       @                ��Ͽk�?wgL����?                                ?���@��?      �?                                                                              �?      @�����9�?��{q��?              �?      �?      �?      �?      �?       @               @       @       @       @       @       @       @              �?c9��?�Y�8��?                                              �?              �?                                                              �?       @�9�፿�?�h�l��x?      �?              �?      �?(�K=�?      �?       @      �?       @       @       @       @       @       @       @              �?��C��?������?              �?                6��9�?      �?              �?       @       @               @       @       @              �?      @e0
84��?��`>�^�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?               @-h#���?���Ű�?      �?      �?      �?                              �?                                                                               @?�]�FR�?�9�:�G?      �?      �?                3~�ԓ��?      �?       @      �?       @       @       @               @       @              �?        x�/���?I����?      �?                         �
���?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?-h#���?���?�?      �?              �?      �?v�'�K�?              �?                                       @       @       @       @                �Po���?�F����?      �?                        �]�����?      �?                       @                       @                                      @xwwwww�?�+�gW;�?                                e�v�'��?              �?               @                       @               @      �?                ��j1v�?�!���\�?      �?              �?        �RO�o��?      �?                       @       @               @                       @      �?      @z�D_r�?�Mܬ�?                              �??���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?        n��W�?����?                                              �?                                                                              �?      @����e�?���W�g?      �?                        �K=��?              �?               @               @       @       @              �?      �?        *L����?0Z���c�?              �?                ���@��?      �?       @      �?       @       @                                              �?       @"�
���?�)��=�?      �?                        �z2~���?      �?              �?                                               @              �?        �`�AQ��?WlϮvD�?      �?              �?      �?��V��?      �?                       @               @               @       @      �?              �?F��s��?��Rî��?              �?                �'�K=�?      �?       @      �?                               @       @       @                       @�������?!N�� �?      �?                        ?���@��?              �?                                               @       @              �?       @�9�፿�?`-��_�?      �?                      �?{2~�ԓ�?              �?               @       @               @                      �?              @s��2�?a�,����?      �?                        !�
���?      �?              �?       @                               @              �?              @�^<���?��l��_�?                      �?      �?F���@��?      �?                                                               @                       @ae��	�?����K#�?      �?      �?      �?        ��ۥ���?      �?       @      �?       @       @       @               @       @              �?       @���-�j�?\)Խ�i�?                      �?        v�'�K�?      �?       @               @       @       @                               @                7O�)��?6��p�?              �?      �?        ���@��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @��Po��?��MP�?                                �@�6�?      �?       @      �?       @       @       @       @       @       @              �?        6��w���?���
��?                      �?      �?F���@��?      �?                       @       @       @               @              �?               @{+�oM�?i�%��?                                ��RO�o�?      �?              �?                       @                                               @k� 6\.�?�����?      �?                        P�o�z2�?      �?       @      �?               @       @       @       @       @      �?               @��l��?��>n�?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?�����%�?                                ?���@��?              �?               @       @                                              �?       @��*��?�c��t"�?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?                       @                              �?      �?        ����+�?�n����?              �?                �K=��?              �?                       @       @               @       @              �?       @��s��2�?͇;Y��?                                ���Vج?      �?              �?               @                       @                      �?      @ J�hY�?���座?                                p�z2~��?      �?       @      �?               @       @               @       @              �?       @�]�FR�?f;=����?                                �@�6�?      �?                       @       @               @       @               @              �?�d�Q���?��6�>�?      �?                                      �?                                                                              �?      @~PT���?B֜�#�h?                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�Y;���?��^}Ν�?      �?                        �ԓ�ۥ�?      �?       @      �?       @               @       @       @       @       @      �?       @��-��?қ]N��?      �?              �?      �?F���@��?      �?              �?       @                                       @                       @
Sb����?l��̿?      �?                        [as �
�?      �?              �?               @                       @       @              �?       @V�;�RG�?�#�����?      �?                        [as �
�?      �?              �?               @               @                              �?       @��I{+�?�~+?^��?      �?                        ���V؜?      �?       @      �?               @       @               @       @                      @_�ti���?Rgض�j�?      �?                        6��9�?      �?       @      �?       @               @                                      �?       @�iŽ�,�?kߤJ�?                                              �?              �?                                                              �?       @D)-��?]v�{x?              �?      �?        SO�o�z�?      �?       @      �?       @               @               @       @      �?      �?        s[ݧ���?��!���?      �?                              �?      �?       @      �?               @       @       @       @       @       @                m�\d���?1�}ܜ�?      �?              �?      �?�RO�o��?      �?                       @       @       @       @                      �?      �?        3���O�?=�k�S��?                                              �?              �?               @       @                                      �?       @]��#�d�?&��=m~?                      �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @                �����`�?���}E��?      �?              �?      �?�]�����?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @b��1��?5OؾI�?                      �?      �?��Vؼ?      �?       @                       @                                              �?      @��W��?���:��?                      �?        ��RO�o�?      �?              �?       @                       @       @       @      �?      �?      �?%���?�4}u��?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�d�Q�ϰ?i�)K�^�?      �?                        �ԓ�ۥ�?      �?       @      �?                                       @                               @S,?(��?Y� ����?      �?      �?      �?        �K=��?      �?              �?                                                                      �?~PT���?��/���?                      �?        �'�K=�?      �?                       @       @               @       @               @      �?      �?3NaJ̖�?���r�R�?                      �?      �?H���@��?      �?       @      �?               @                       @       @      �?              @
�R,�?�Yk��-�?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                      @Y�)L�ْ?)�<$3�?      �?                              �?              �?               @               @       @       @       @       @      �?      �?q���Y�?���X$�?      �?              �?      �?��V��?      �?       @               @       @       @                       @      �?              �?7��`�A�?#�$g��?      �?              �?      �?��RO�o�?      �?       @      �?       @       @               @       @                               @��¯�D�?4!F1�}�?      �?              �?        ?���@��?      �?              �?                                       @                      �?       @���!���?H���?                      �?              �?      �?       @      �?               @       @               @       @      �?      �?       @�^<��u�?f̮����?      �?              �?              �?      �?       @      �?               @       @       @       @       @       @      �?      �?��"s�g�?��w�T�?      �?              �?        �@�6�?      �?       @      �?                       @       @       @       @              �?       @)����?W)5M:z�?      �?              �?      �?6���?      �?       @      �?                       @       @               @       @                |]�;�?��8�y�?      �?              �?        ��V��?      �?                                                                              �?      �?�9�፿�?�SQS�?                      �?        F���@��?      �?                                                                      �?               @�vAIE�?ƸI��?                                              �?              �?                                               @              �?       @9�WH�?����}?                      �?      �?Zas �
�?      �?       @               @       @       @       @               @      �?      �?       @)�tN|x�?=k��?      �?                        �@�6�?      �?                                                                                      �?���8�)�?R9���?              �?                �6��?      �?                       @       @                                              �?      �?�i����?�6.�{�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @                ^��Z��?L@��Z�?      �?                        �D+l$�?      �?                       @       @               @       @              �?               @�V�ߚ�? �����?      �?                        H���@��?      �?              �?                       @       @       @       @       @                ��E���?-?�Hl�?                                F���@��?              �?                               @               @       @                       @���w��?m��ݠ�?      �?                        SO�o�z�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @?�]�FR�?--����?                                ��Vؼ?      �?              �?                       @                       @              �?      �? J�hY�?]f(���?      �?              �?        F���@��?      �?       @      �?                       @               @       @              �?      �?{�rv��? U\:���?                      �?        3~�ԓ��?      �?       @      �?               @       @       @       @       @              �?       @���(���?L��N�?      �?              �?      �?�6��?      �?       @      �?                       @               @       @              �?      �?�3i�ae�?�5vl�?      �?              �?      �?�K=��?              �?               @                                              �?                ���J�?��L,�?      �?                        �'�K=�?      �?              �?                       @       @       @       @              �?       @�^<��u�?�N>���?                      �?              �?      �?       @               @       @       @       @       @       @       @                :Blӊ{�?�#M���?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?        E�Ή�?;���P
�?      �?              �?      �?�V�H�?      �?                       @               @       @       @       @       @              @�����?�]t�dD�?      �?              �?      �?      �?      �?              �?       @       @       @       @       @       @       @                WH�%���?�H���?                                              �?       @       @      �?      �?      �?      �?      �?      �?              �?      @�rv��?���,�GJ?      �?              �?        ��ۥ���?      �?       @               @       @               @                       @                �������?=�u#�7�?                              �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?                      �?n��W�?�@�ª?              �?                �]�����?      �?              �?       @       @               @       @       @              �?      �?kH����?��9I��?      �?              �?      �?�@�6�?      �?              �?                                       @                      �?        �?^���?C���?      �?              �?      �?      �?              �?               @       @       @       @       @       @       @      �?      �?��M+��?�x��x�?                                              �?               @      �?      �?      �?      �?      �?      �?                      �?�'�F7�?O���&?      �?                                      �?              �?                                                              �?       @�bѲ
n�?�9.�� x?      �?              �?      �?�@�6�?      �?                               @       @                                      �?      @��W��?	s���?      �?                              �?      �?       @               @               @       @       @       @       @              �?�H*���?%Y��N�?                      �?      �?ܥ���.�?              �?                                       @                              �?      �?�1���? �d	Ž�?      �?              �?      �?��RO�o�?      �?                       @       @               @       @               @      �?      @K��a�?��h�g�?                                ?���@��?      �?              �?       @               @       @               @              �?        �FR,?�?RMM2�å?                      �?        ���Vج?      �?              �?                                                                       @��j1v�?�b��e�?                      �?        p�z2~��?      �?              �?               @       @               @       @              �?      �?��E���?��u/��?                                �'�K=�?      �?                               @               @       @                      �?       @_W-��?)H���?                                              �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?@Ր�,?                      �?      �?6���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?qi��|��?3��+�?                              �?�@�6�?      �?       @      �?               @                       @                      �?        ��|�?^�?�C���?      �?                      �?>�]���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�r@��?O�9��?      �?              �?              �?      �?       @                       @       @       @       @       @       @      �?        Ͽk�.M�?,"4D�@�?                      �?        ���V،?      �?              �?                                                              �?      �?�V�ߚ�?�F����?      �?              �?      �?v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @E�(Ţe�?��-9y��?      �?              �?        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?E�(Ţe�?B�s�[��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�U�����?qpTV�?      �?                        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        nC��x�?A{��d�?      �?                        �@�6�?      �?              �?               @                       @                      �?       @��>|]�?n��k�Ϋ?      �?                        6��9�?      �?       @               @       @       @       @                      �?               @�����T�?��#����?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?                               @       @       @       @      �?       @E������?���?�?      �?                        Zas �
�?              �?               @       @       @       @       @               @              @؋�ߵN�?ltB%��?      �?                        �'�K=�?      �?       @      �?                                               @                        �s��2�?��n��?                                SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        nC��x�?nm�'�c�?      �?      �?                �@�6�?      �?                                                                                      �?f��	��?����Ys�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�U�����?~s���+�?      �?      �?                p�z2~��?      �?       @      �?                                       @                      �?      �?�����?"L�q�h�?      �?      �?                [as �
�?      �?       @      �?               @                       @                      �?       @j��|��?���Z���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @Y�)L�ْ?3<�O��#?                      �?        (�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                ����'t�?$������?                      �?        ��ۥ���?      �?       @      �?       @       @       @       @               @       @      �?      �?g�����?Ih���-�?                                �K=��?      �?       @      �?       @       @       @               @                      �?      �?%��}��?E~�[�?                      �?        SO�o�z�?      �?       @               @       @               @                              �?      �?�w�ӥ��?�P�~��?                      �?        Zas �
�?      �?       @      �?       @       @       @                                               @j��|��?��G��?              �?      �?        ܥ���.�?      �?       @      �?       @       @       @       @       @       @                       @/h#���?��찣�?                                F���@��?      �?                       @                       @                      �?              @�a/��?�� ;�c�?      �?                        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @^��Z��?�~�θ�?                                p�z2~��?      �?                                       @       @       @       @       @              @�@ʾ���?�RW���?      �?      �?      �?        ,l$Za�?      �?       @      �?               @                               @      �?              @Z;��V�?Cbm6��?                      �?        H���@��?              �?                       @               @       @       @      �?      �?      �?|]�;�?֪�sze�?                                �ԓ�ۥ�?              �?               @       @               @                      �?      �?      @h�����?�6��y�?                              �?��RO�o�?      �?       @      �?       @                       @                              �?      @�6��w��?�[zmo��?      �?              �?      �?      �?              �?               @       @       @                               @              �?����?p7,"4D�?      �?                        v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?       @                ^��Z��?! `��=�?                      �?      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �bѲ
n�?x��u�v�?      �?      �?      �?        e�v�'��?      �?       @      �?                                                                        �/�Q��?�ơe��?      �?                        ?���@��?      �?       @      �?                                                              �?       @,�����?r���"�?              �?      �?        �RO�o��?      �?              �?       @       @       @       @       @       @       @      �?        �d�#�6�?���׍�?                      �?        ��.�d��?      �?                       @               @               @              �?      �?      @��Z�KS�?|Y���?      �?                        ��.�d��?      �?              �?               @       @       @       @       @      �?      �?        e0
84��?��q�?��?      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @               @�፿Po�?(h����?      �?      �?      �?      �?      �?              �?               @       @       @       @       @       @       @      �?        1�z�Τ�?��8�g�?                                �'�K=�?      �?                       @       @       @       @       @       @                      @#���?�xN����?      �?                        �
��V�?      �?       @                               @               @       @       @      �?        �Q����?1>�T6��?      �?                        ��.�d��?      �?              �?       @               @               @              �?               @�`ph>�?�n�\m�?      �?                        ���@��?      �?              �?       @       @       @       @                      �?      �?      �?C)-���?Ʌ�ֺ�?                                �'�K=�?      �?                                                       @              �?              @z����"�?�"ѽ@��?      �?                        �ԓ�ۥ�?      �?       @               @               @               @                              @>�/�Q�?����p�?      �?                      �?F���@��?      �?              �?                                       @                      �?      �?c=kg��?5�F����?      �?              �?        ��.�d��?      �?       @      �?               @               @               @              �?      �?�:��?2��O��?                                �o�z2~�?      �?       @                       @       @       @       @       @       @                �s��2�?~C��`�?      �?                        $Zas �?              �?               @       @               @       @                      �?      �?��<݌�?���5π�?      �?              �?        �z2~���?      �?              �?       @       @       @                                      �?       @l	�Y �?�uy9 ͻ?      �?                        �o�z2~�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?n��W�?�_k�x�?                                �]�����?      �?       @      �?                                                      �?      �?      �?T�n�Wc�?���?                                              �?              �?                                                                       @}�?^��?ľl�ox?              �?                      �?      �?       @      �?               @       @       @       @       @       @      �?        �KS}��?�����?      �?              �?      �?�]�����?      �?                                               @                              �?       @��x�]��?N�����?                                ,l$Za�?      �?              �?               @       @               @                      �?      �?�E�*�A�?��X74�?      �?      �?      �?        H���@��?      �?       @      �?               @                               @                      �?�^!ї��?���r¸�?      �?              �?      �?�o�z2~�?      �?                       @               @       @               @      �?              �?5�u�b��?	����?              �?                �ԓ�ۥ�?      �?                               @                                              �?      �?h#���?%y���?                      �?      �?�@�6�?      �?              �?                       @               @       @              �?        p2��g�?�� �G�?      �?                                      �?              �?                                                              �?       @�vAIE�?�!��}�w?      �?                                      �?                                       @       @                                      @�፿Po�?\��J5"q?      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @ś�8j��?JޣT�0�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�U�����?tq]�?      �?                        �K=��?      �?                       @               @                       @       @                �*��?�S=z7	�?                                p�z2~��?      �?       @      �?               @       @               @       @              �?       @q���Y�?�����H�?                      �?        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                        nC��x�?��*�!�?                      �?              �?      �?       @      �?       @       @       @       @                       @      �?        rv��?&E�r�)�?      �?              �?      �?p�z2~��?      �?       @               @                       @       @       @                        �����?:$F�f#�?      �?                        6��9�?      �?       @               @       @       @       @       @       @      �?      �?        ���l	�?�h��W��?                      �?      �?�
��V�?      �?              �?       @                                       @      �?      �?        �Po���?��_- �?                      �?      �?�ԓ�ۥ�?      �?                               @       @       @                      �?                i1v��?D�!��e�?                      �?      �?�RO�o��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?]����`�?`�Ö��?      �?      �?                ���Vج?      �?              �?                                                              �?      @��w����?mt���?                                �]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @]����`�?V�uiC�?                      �?        �o�z2~�?      �?       @      �?       @       @       @       @       @       @       @              @��3��x�?�\�V�`�?                      �?      �?�K=��?              �?               @       @       @       @       @               @              �?�
����? ����?      �?      �?                              �?              �?                               @                                       @�6��`��?5� ��kz?              �?                Zas �
�?      �?       @      �?                                       @       @              �?       @M��o2��?�6����?      �?                        �V�H�?              �?                               @       @                      �?              �?���w��?�}`�o�?      �?              �?              �?      �?       @                       @       @       @       @       @       @      �?      �?b�(Ţe�?{5��?                                ��.�d��?      �?                                       @                       @              �?       @H���<�?�J��V�?      �?              �?      �?�'�K=�?      �?       @                       @       @               @       @                      �?���U���?�ӯ�2�?      �?                        F���@��?      �?       @      �?       @                               @       @                      @��	�p�?�V�j���?      �?              �?        �z2~���?      �?       @      �?               @       @                                               @~5&��?�%�g���?      �?                      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?                      �?����[�?��'q�?                      �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�X����?�c����?      �?              �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�Y;���?�[�N�ɰ?                      �?              �?      �?       @               @       @       @               @       @       @      �?      �?�%��f��?o�w{���?                      �?      �?SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @m+�oM�?���C�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?9�%��}�?�����?                      �?        ��ۥ���?      �?       @               @       @       @       @       @       @       @              �?}�mu��?S���p��?      �?              �?      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?               @�X����?BAM�<.�?      �?      �?      �?        6��9�?      �?       @      �?                                       @       @              �?       @�-�jL��?��WtJ��?                      �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @^��Z��?nWʜKa�?                      �?        �K=��?      �?       @               @       @               @                                       @��>�MF�?����e��?                      �?              �?      �?       @      �?       @                                               @                *L����?RY�f �?              �?                ��ۥ���?      �?       @               @       @       @       @       @       @       @              @t3NaJ��?�	��r+�?                      �?      �?���Vج?              �?                                                                              @?�]�FR�?%s�I7�?      �?                        �'�K=�?      �?       @                                                                               @;��u�4�?���i��?                      �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        Rp�l?�X��ep�?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @����'t�?g�`F<3�?              �?      �?        �D+l$�?      �?       @      �?       @       @       @       @                      �?      �?       @z����"�?=�V�-.�?                      �?      �?	��V��?      �?       @                               @       @                      �?      �?      @M|x�/��?ʉ����?                                6��9�?      �?       @      �?       @       @       @                                                	�U:�?��y��?                                �'�K=�?              �?               @               @       @                      �?      �?      �?H���<�?���v��?      �?                        ���.�d�?      �?       @      �?       @               @       @               @       @              �?����?Mhe:r�?                      �?      �?��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?       @              @E�(Ţe�?
'�y\�?      �?              �?      �?�z2~���?      �?                                                       @                      �?      @|]�;�?$#"W��?              �?                ��RO�o�?      �?              �?               @                                              �?      �?��[��?;Y�)n�?      �?              �?      �?�]�����?      �?       @      �?                       @       @       @       @      �?      �?      �?��0%f�?�.}ޓ^�?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @              �?���9���?]Ӂ�wX�?      �?                        ���@��?              �?               @                       @                      �?      �?      @�������?8H ����?                      �?        6���?      �?                       @       @                       @                      �?      �?��M+��?{&����?      �?      �?      �?        ��V��?      �?              �?                                                      �?      �?        Y�ڙ���?�נTF��?                      �?        p�z2~��?      �?       @      �?                       @                                      �?      @��<݌�?2����5�?              �?      �?      �?��ۥ���?      �?       @               @       @                       @              �?               @�c9�?K���3T�?                      �?      �?��V��?      �?       @               @       @       @       @       @       @       @                ^!ї�V�?pQ����?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @-h#���?"�O4�?      �?              �?        SO�o�z�?      �?       @      �?                       @       @       @       @      �?      �?       @�v&�1��?��(���?      �?                        �D+l$�?      �?              �?               @                       @       @      �?      �?        rv��?gi($�,�?                      �?              �?      �?       @               @               @       @       @       @       @      �?         ʣ��8�?����S�?      �?              �?      �?�]�����?      �?       @               @                       @               @      �?      �?      �?��m$�?�찣L�?                                      �?      �?       @               @       @                                       @                <�RG�m�?��]3�[�?                                              �?               @      �?      �?      �?      �?      �?      �?                       @�Y;���?��ֺ�,?              �?                �@�6�?      �?              �?                                       @       @              �?       @�G�Ɉ��?�U$��7�?                                ���V؜?              �?                                                                               @��N�Ա?� ��r?                      �?        ���@��?      �?       @      �?       @       @               @       @       @      �?               @�l��?���
��?                                �ԓ�ۥ�?      �?              �?               @       @                                               @�Q����?S!��?      �?              �?        (�K=�?      �?              �?       @       @       @       @               @       @              �?mӊ{'Y�?�7J-�?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?�q0|��u?                                ��RO�o�?      �?       @      �?       @       @       @                                               @�?y4��?�c|A�?      �?                        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                ����'t�?/ɾ.Y�?      �?                        p�z2~��?      �?              �?               @       @       @                              �?       @l�\d��?_}���?      �?                        ���V،?      �?                                                                                      @ui��|��?Ѯ^� f}?                                �'�K=�?      �?       @      �?                                                              �?      �?����9��?o%��Q�?      �?              �?        ��Vؼ?              �?                                       @       @                              @�U�����?6��X�R�?      �?              �?      �?�]�����?      �?                       @               @       @       @              �?      �?        �Q���\�?،p�K��?      �?              �?      �?      �?      �?       @               @               @       @       @       @       @      �?      �?kg����?��>n�?      �?                        H���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @����[�?Q�.}ޓ�?      �?      �?                Zas �
�?      �?       @      �?                                       @                      �?       @�&`��?����?                      �?      �?�'�K=�?      �?       @      �?               @       @               @       @              �?        �������?�<a���?                                �'�K=�?              �?                                                                      �?      �?\��r�?O\����?      �?      �?                ���Vج?      �?              �?               @                               @              �?       @�}�m�?�d�(�?                      �?        6��9�?      �?       @                       @               @               @      �?              @���q%�?�_7r~�?      �?                        ���Vج?      �?       @                                                                               @�c=kg�?��N�%�?                      �?      �?�@�6�?      �?                               @                       @              �?      �?      �?�E�X���?��4'ʬ�?      �?      �?                �@�6�?      �?              �?                                               @              �?      �?Y���d�?�w?�?      �?                        p�z2~��?      �?       @               @                                                      �?        ;�^!��?�8�>�h�?      �?                                      �?                                                                                      @X�ڙ���?x c[�ch?                      �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?F��1��?��-wZ�?                      �?        {2~�ԓ�?      �?       @                       @                       @              �?                �C��?��k�4R�?      �?              �?      �?�
��V�?      �?                       @                                       @      �?              �?H���<�?kZ�P-�?                                6��9�?      �?              �?       @               @       @       @       @              �?       @Ɉ���!�?� �{K�?      �?              �?        ��V��?      �?       @      �?               @       @                       @              �?       @Τ=����?j�j�6��?                                6��9�?      �?       @               @                               @              �?                ���Z��?>K sQ3�?                      �?      �?H���@��?      �?       @      �?                       @                       @              �?       @R��'��?�-�+Z�?                      �?              �?      �?       @      �?       @       @                                       @      �?        
Sb����?Oʿ�pG�?      �?              �?        ,l$Za�?      �?                       @       @               @                      �?      �?        G�%��}�?�.骀�?      �?                        P�o�z2�?      �?       @      �?       @       @       @                       @       @      �?        1@�bѲ�?�2Ĥ�T�?      �?              �?        �ԓ�ۥ�?      �?       @      �?       @                               @       @              �?       @	{�����?�e�Haw�?                                ���V؜?      �?                       @       @                                                       @c9��?h[�ɎL�?                      �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?        8�]�FR�?��R���?      �?              �?        (�K=�?      �?       @               @               @       @               @       @      �?      �?	�{B��?�ct�E��?      �?                        ���V،?      �?              �?                                               @              �?       @ZV����?氾6�-�?      �?              �?        H���@��?      �?       @               @               @       @       @       @      �?               @����?7{Č��?      �?                        �ԓ�ۥ�?      �?       @      �?               @                                              �?       @7w\I`��?����*�?      �?              �?        �ԓ�ۥ�?      �?       @      �?       @       @       @       @       @       @       @      �?        }�mu��?Pm���?                      �?        �ԓ�ۥ�?      �?              �?                       @               @       @              �?      �?q��3���? ����?      �?                        ���V؜?      �?       @                                       @       @                      �?      @��M+��?l8sI���?                                $Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�Y;���?1{�����?              �?      �?      �?�
��V�?              �?                                               @                      �?       @3\.2�z�?J|��4�?      �?                        ���V؜?      �?                                               @       @       @              �?       @�vAIE�?*�t�c�?                      �?      �?!�
���?      �?              �?       @       @                                              �?        Y���d�?�)ǉ��?                      �?        H���@��?      �?       @                                                                      �?      �?�����?���O��?      �?                                      �?              �?                                                              �?       @%�yO�0�?#��=�w?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?              �?       @n��W�?:yl����?      �?      �?      �?        ���V،?      �?              �?                       @               @       @              �?      �?��[�՘�?��_*>�?                      �?        �'�K=�?      �?       @      �?                                               @              �?      �?��`�AQ�?m�
]~��?      �?                        $Zas �?      �?                                               @                       @      �?        ፿Po�?|P��@��?                                $Zas �?      �?                                                                              �?       @��J��?�D�Tպ?                                �z2~���?      �?       @      �?                       @                       @              �?      �?}�mu��?~#*��?      �?      �?      �?        3~�ԓ��?      �?       @      �?               @       @               @       @                        ����>�?ˢ���?      �?              �?        Zas �
�?      �?       @      �?               @               @       @               @      �?       @=���&�?��"��?                      �?        !�
���?              �?                       @                       @       @              �?       @O�)���?#M�ַ�?                      �?      �?��RO�o�?              �?               @       @       @                       @              �?        Y���d�?w�i+�I�?      �?              �?      �?�6��?      �?       @               @               @       @       @       @       @      �?        ��3i�a�?��.��5�?      �?                        ��Vؼ?      �?                       @               @       @       @                      �?      @>�/�Q�?gv|���?                      �?      �?��RO�o�?      �?       @       @      �?      �?      �?      �?      �?      �?                      @<݌S��?7�����?              �?                H���@��?      �?       @      �?       @       @       @       @               @      �?                ���-��?������?                                              �?                       @                                                      �?        ���Y;�?ϾGH;l?      �?                                      �?              �?                                                              �?      @~PT���? ��j��x?      �?                        �z2~���?      �?              �?       @       @       @       @       @       @      �?              �?&>����?�чڂ�?                                ���Vج?      �?       @      �?                                       @       @              �?      @1[�yj�?�fQ0��?              �?      �?        p�z2~��?      �?       @      �?       @                                                               @���!���?Ŏ����?      �?                        ��ۥ���?      �?                               @               @               @      �?      �?      @}�mu��?��n��O�?              �?      �?        >�]���?      �?       @      �?                               @                              �?        HE�����?���&8p�?                      �?      �?�]�����?      �?                               @                       @       @      �?      �?        >�/�Q�?R������?      �?              �?        ��RO�o�?      �?       @      �?                                               @              �?       @Ͽk�.M�?�g�x��?                      �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?                      @#w\I`ޓ?�/�a_x�?                      �?      �?e�v�'��?      �?       @               @       @       @       @       @       @       @              �?�+	�{B�?����C�?                                ��Vؼ?      �?              �?                                       @                      �?        {������?�È��?      �?      �?      �?      �?��.�d��?      �?       @                       @       @               @       @      �?      �?       @B�/����?�ֲAH��?      �?      �?      �?        3~�ԓ��?              �?               @                       @                      �?                f{����?K�*����?      �?      �?                �K=��?      �?              �?                                                                      �?�Kn��4�?���Ʃ�?                      �?      �?>�]���?      �?       @               @               @                       @      �?      �?        ����`�?1�^O���?                                ���V؜?      �?       @      �?                                                                        �u�b���?��s1G�?              �?      �?      �?      �?      �?       @               @       @       @       @       @       @       @      �?        �
����?���O��?      �?      �?      �?        �D+l$�?      �?       @      �?                                                                      @K�ć7��?M�E�:�?                                ��Vؼ?      �?              �?       @                                                      �?      �?��N���?�C$#"W�?                      �?      �?��RO�o�?      �?       @       @      �?      �?      �?      �?      �?      �?       @               @Xph>ׯ?�y���?      �?              �?      �?P�o�z2�?      �?       @                       @               @               @       @              �?o��z��?pؓ [��?                      �?        !�
���?      �?              �?                                                                      @�Kn��4�?���pj��?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�U����|?�ᦵ�?      �?                        3~�ԓ��?      �?              �?       @       @       @       @       @       @       @              �?m�\d���?�Zi�a��?      �?                                      �?       @      �?               @                                              �?       @Y���d�?����G�|?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?Rp�l?��*,M�?                      �?        P�o�z2�?      �?       @      �?       @       @       @               @       @       @      �?        ����w�?���5���?                      �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?��1�~?���m��?      �?              �?      �?$Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @              @n��W�?�2�R���?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                h��2�?$�E���?                      �?        �'�K=�?      �?              �?       @               @               @       @                       @۴��I��?�R�Ea�?                      �?              �?      �?       @               @               @       @       @       @       @      �?      �?a�:�?	F9q�?              �?                �
��V�?      �?       @      �?                       @       @       @       @              �?       @{B���?P�$�5�?                                ���V؜?      �?       @      �?                                                                       @�cX�~k�?�8n��7�?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              @F��1��?�2�*.�?      �?      �?      �?        	��V��?      �?              �?                                               @                        +�d�#�?��b�Z�?              �?                ���V،?      �?              �?                                                              �?       @�r@��?)ε&�2�?                      �?        ���.�d�?              �?               @               @       @               @       @               @o�)L���?f�[$�?      �?                        $Zas �?      �?       @                                       @                       @      �?      �?[ݧ����?�$g��?                                 �
���?      �?              �?                                                              �?      �?b����,�?��`6F��?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?�Ѱ{�?                              �?	��V��?      �?                                                       @       @              �?      @&��f���?V2�P��?                                              �?               @      �?      �?      �?      �?      �?      �?                      �?-h#���?��??      �?                        �z2~���?      �?                               @               @                              �?      @N��b��?5^��1��?                                �]�����?              �?                               @               @       @              �?        ��*��?5xc�?                      �?      �?e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        E�(Ţe�?%������?      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?       @                E�(Ţe�?�����?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @m+�oM�?�
�!��?      �?              �?      �?�K=��?      �?                       @               @       @                       @      �?        a/���?��pY�?                      �?        ��RO�o�?      �?              �?       @       @       @       @       @       @      �?               @=P9��_�?E����z�?      �?      �?                �'�K=�?              �?                               @                                      �?       @�����f�?HƓf���?                      �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @                m+�oM�?�1RT P�?                      �?         �
���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @!�iŽ�?/-��禳?      �?                        ��RO�o�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ���Z��?�������?      �?      �?      �?        H���@��?      �?       @      �?       @                                       @      �?      �?       @B����?�g�EQ��?      �?              �?        �z2~���?      �?       @      �?               @                                                        �X����?�i����?      �?              �?                              �?                                                                      �?       @9�%��}�?�5(�A?      �?                        �'�K=�?      �?       @      �?                                       @              �?      �?       @}x�/���?RoS�Q+�?      �?                        �6��?      �?                                       @       @               @      �?      �?      @����>�?-��7u@�?      �?                        ��RO�o�?              �?                       @                                              �?      @�7�B�]�?T����?                                p�z2~��?              �?               @               @       @                       @              @�*��?�Tv�k�?              �?                ���V؜?      �?                                                                                       @�{'Y��?�eXg��?                      �?      �?	��V��?      �?              �?                       @       @       @       @      �?                �Τ=���?�-d����?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @Y�)L�ْ?3<�O��#?              �?      �?        �D+l$�?      �?       @      �?               @                       @                      �?       @�^!ї��?�p�uC�?                      �?        �'�K=�?      �?              �?               @                                                        k� 6\.�?w�u�C/�?      �?              �?        Zas �
�?      �?       @      �?                                       @       @      �?      �?        ӊ{'Y��?�TͿ���?      �?              �?        ?���@��?      �?              �?                       @       @                              �?      @r�g�L��?�!����?                                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�%��}�?� �?      �?              �?      �?�K=��?      �?       @      �?               @       @                              �?               @dsǕ�?��1bJ��?              �?      �?                      �?               @      �?      �?      �?      �?      �?      �?              �?      @9�%��}�?��8�/?      �?                        �ԓ�ۥ�?      �?                       @                                                               @��r�9��?��2pI�?      �?              �?      �?              �?                                                                                       @�9�፿�?��Y�pWh?      �?              �?        �RO�o��?      �?               @      �?      �?      �?      �?      �?      �?       @              @8�]�FR�?^3�[?N�?      �?                        ���V،?      �?              �?               @                       @       @                       @�:��?��r��?                                �]�����?      �?       @               @                       @                              �?      @䛌8j��?J9�3�<�?              �?      �?        $Zas �?      �?                               @                               @              �?       @ٴ��I��?�Ψ��R�?                                [as �
�?              �?               @       @               @               @       @      �?        h#���?��p��,�?      �?              �?        �]�����?      �?               @      �?      �?      �?      �?      �?      �?              �?        1[�yj�?�r#Hǿ�?      �?              �?      �?��RO�o�?      �?       @                               @       @       @       @      �?      �?      @?^��C�?I�L}��?      �?              �?      �?$Zas �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @��>�MF�?X6��$�?      �?      �?                �'�K=�?      �?                                       @       @                      �?      �?       @��Dz�r�?4�G�?              �?                ��.�d��?      �?       @      �?       @       @       @               @       @                      �?�KS}��?F�)�#~�?      �?              �?      �?3~�ԓ��?      �?              �?       @       @                               @      �?      �?       @�?y4��?|>XT^1�?                      �?      �?(�K=�?      �?       @      �?       @       @       @       @                       @                1[�yj�?o�\m9�?      �?                        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                3�$0�	�?�T�?      �?              �?        �ԓ�ۥ�?      �?       @      �?                                       @       @              �?       @&���[�?��ZY��?      �?              �?      �?      �?      �?       @      �?               @       @       @       @       @       @      �?        ��M+��?��./��?      �?      �?      �?        �'�K=�?      �?       @      �?               @       @                       @              �?       @�	�p��?w�"�?                      �?        P�o�z2�?      �?       @               @       @       @       @                       @              �?��=���?8x���?                                ���V،?              �?                                                                               @Xph>ׯ?d��"j?      �?                        �K=��?      �?       @      �?               @               @       @       @              �?       @�������?Z��$o�?      �?                        ���@��?      �?              �?       @       @               @               @              �?      �?����?�X�|v�?                                ���V،?      �?              �?                                               @                       @��r�9��?]��F��?                      �?        �@�6�?      �?                                               @                              �?       @���w��?���c�Ɲ?      �?                        ���V؜?      �?              �?                       @       @       @                      �?      @t3NaJ��?�r�ة�?                      �?        ��ۥ���?      �?                       @       @       @       @       @       @      �?      �?        y4��0�?=+���A�?                      �?      �?      �?      �?       @      �?               @       @       @               @       @      �?        �������?y>��A�?      �?                        6��9�?              �?               @       @               @                       @      �?      @�����f�?��D�?                                �ԓ�ۥ�?      �?              �?                                                              �?       @�/�����?��EA�&�?      �?      �?                p�z2~��?      �?       @                       @                                                      �?R��'�F�?���@���?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?                       @]����`�? <���9?      �?                        ���Vج?      �?                               @                                              �?       @$���?@=_�Ŝ?                                ��RO�o�?      �?                       @                                                                9�WH�?�+�r^g�?      �?      �?      �?        H���@��?      �?       @      �?       @       @       @                                      �?       @M���E�?���|W��?                              �?              �?                       @                                                              @���'�?Ѯ^� fm?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�%��}�?țmͷ�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @����[�?wWVU�%�?      �?              �?      �??���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?nC��x�?��)��q�?      �?      �?      �?        Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                )g��1�?�g�Y��?      �?                        {2~�ԓ�?              �?                       @               @                      �?              �?L��b��?�+5�%�?      �?              �?      �?P�o�z2�?              �?               @       @       @       @               @       @      �?      @�0%fK�?��5vl�?                      �?        ��ۥ���?              �?                       @       @       @       @       @       @                �C��x�?V��Y�z�?                      �?        �K=��?      �?       @      �?                       @               @       @              �?       @
�R,�?K�ù7�?                                �6��?      �?               @      �?      �?      �?      �?      �?      �?       @              @n��W�?�X�]Y�?      �?                        �z2~���?              �?                       @               @                                      @Y�՘H�?(��?                                {2~�ԓ�?      �?       @      �?                                               @                        �'�F7��?�O4����?                      �?        �]�����?      �?                       @               @       @       @       @       @      �?       @)���G�?�-l�j�?      �?              �?      �?$Zas �?      �?                       @       @       @                              �?               @�^<��u�?IH�w�+�?                      �?        P�o�z2�?      �?                       @                       @                      �?                ������?�\RI�?              �?                ��ۥ���?      �?       @      �?       @       @               @       @              �?      �?      �?�p����?3+�^�r�?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @�፿Po�?�V�φn?      �?              �?              �?      �?       @      �?       @       @               @               @       @      �?        ���?y4�?�C��?                              �?Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?)g��1�?�/׽~��?      �?              �?      �?�o�z2~�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �r@��?N�D%��?      �?              �?      �?�@�6�?      �?                                                                              �?        X�ڙ���?�+� n��?      �?      �?      �?        �'�K=�?      �?       @      �?                               @                              �?       @���Up�?N��k��?                      �?      �?���V،?              �?                                       @                                        
�X����?��ׇh?      �?                      �?��ۥ���?      �?       @      �?       @               @               @       @       @                Q�n�)�?l5��0�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @����'t�?&����?                                ���V،?      �?                               @                                                      @��̱���?s	�f�?      �?              �?      �?!�
���?      �?       @      �?       @       @               @       @       @      �?              �?b/��:�?����?                                ���V،?      �?                               @               @                              �?      �?�፿Po�?kYE3�փ?                      �?              �?      �?       @               @       @       @       @       @       @       @                ��r�9�?����\�?                      �?      �?3~�ԓ��?      �?       @      �?       @                               @                               @�=����?&�\��J�?      �?                        v�'�K�?      �?              �?       @               @       @       @       @       @      �?        O|x�/��?���[4�?      �?      �?      �?        (�K=�?      �?              �?       @       @       @               @       @       @              �?�������?�*�@��?      �?              �?        �D+l$�?      �?       @      �?                                               @      �?               @�}�m�?ϱ8Ĵ�?                      �?      �?�@�6�?      �?                       @                       @       @       @      �?      �?      �?�6��`��?�j��g�?              �?                ���V؜?      �?              �?                       @                                              @��C��?�������?      �?                      �?�6��?      �?       @      �?                       @               @       @              �?        ����?^l���?      �?                        ���V،?      �?              �?                                                              �?      �?�Z�<��?�6͉2k�?                                �@�6�?              �?                       @                               @              �?       @�S��%�?߸�9��?      �?                        [as �
�?      �?       @      �?               @                                              �?       @�b��!�?60�\�?                                �z2~���?      �?       @      �?       @                               @                      �?        �^!ї��?i�$d��?      �?                        F���@��?      �?                               @               @       @       @                      @����U��?T�%���?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�m��W�?G��3��?                                (�K=�?              �?               @       @       @       @                       @      �?        X�ڙ���?�_7r�?                                6��9�?      �?                                               @               @              �?      @��8�)1�?.�G��
�?                      �?      �?���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @�j1v�?r2s�I�?                                              �?                               @                                                       @�F���?n�CTm?                                              �?              �?                                               @              �?       @�j1v��?|��h��|?                      �?        �z2~���?              �?                               @               @       @              �?        h#���?,}����?      �?      �?      �?        ��ۥ���?      �?       @      �?               @                       @       @              �?       @ӊ{'Y��?��7m�<�?      �?              �?      �?      �?      �?              �?       @               @       @       @       @       @      �?      �?ߚ ���?~p�L��?      �?      �?                6��9�?      �?              �?                                               @              �?       @�I�:Bl�?�p!���?      �?      �?                6��9�?      �?       @      �?                       @                                      �?       @��*��?�;�/�u�?                      �?      �?�K=��?              �?               @               @       @       @       @      �?              @�N��b�?w�.��)�?                      �?      �?�z2~���?              �?                       @       @       @               @      �?                w�����?J7o���?      �?              �?        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�፿Po�?�:7�6�?                                �D+l$�?      �?       @      �?       @       @       @                       @              �?        �E�X���?v�W�T��?      �?      �?      �?        �K=��?      �?       @      �?                                                              �?       @x�ӥ�>�?�װJ���?              �?      �?        P�o�z2�?      �?                               @       @       @                      �?      �?        �L�5A �?��"R9�?      �?                        ?���@��?      �?              �?                       @                                      �?        	�{B��?�1�X�?      �?                      �?���V؜?      �?              �?                                                                       @�7�B�]�?�}hUDɗ?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?        B6w\I`�?�i%�?      �?                        ��RO�o�?      �?                       @               @       @       @       @      �?               @8q��3�?��߄3�?      �?                        �'�K=�?      �?                               @               @       @                      �?       @�c=kg��?�c�A�?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @E�(Ţe�?�G�O���?                      �?        ��V��?      �?       @      �?               @       @       @       @       @      �?      �?      �?�^!ї�?�P[п7�?              �?      �?        ���Vج?      �?              �?                                                                       @���"X~�?R&�oĠ?      �?                        �
��V�?      �?              �?                       @       @               @                       @�jL�*�?��z]yA�?              �?      �?        (�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�%��}�?�:�<Q�?      �?                      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @-h#���?��N�c�?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @               @ �&#���?1Ȓ:��?      �?              �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @ś�8j��?vV���?                      �?      �?(�K=�?      �?       @               @                                       @      �?                dsǕ��?��%B��?                                �@�6�?      �?                       @               @       @                      �?      �?       @z�rv��?C�� O�?      �?                         �
���?      �?       @               @       @                                      �?               @�+$���?xŚ�?      �?              �?      �?��V��?      �?       @      �?       @               @       @       @       @       @                	�p���?�W�T���?              �?      �?        e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�U����|?2{%r�?      �?              �?              �?      �?       @      �?       @       @       @               @       @       @      �?       @H���<�?Pm��t�?      �?              �?      �?�'�K=�?      �?       @               @       @               @               @       @      �?      �?�.M��o�?2<yl���?                      �?      �?�@�6�?              �?               @                                                      �?       @$X~PT�?�\���[�?                      �?        !�
���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�6��w�?H���?                      �?      �?P�o�z2�?      �?       @      �?               @               @                      �?      �?        �������?^1��?      �?                      �?P�o�z2�?      �?       @               @       @               @       @       @       @      �?        c"=P9��?�k�]6��?      �?                      �?�@�6�?      �?       @      �?                       @                                      �?      @�|�?^�?��Ϟ���?      �?                        ���V،?              �?                               @               @       @              �?       @!�iŽ�?�Ի�?                                ?���@��?      �?              �?                                                              �?        ��=���?i��z	�?                      �?      �?���.�d�?      �?       @                       @                                      �?      �?        [ݧ����?*T�<��?                                �
��V�?      �?       @      �?                                                              �?       @���v�?��Z�x�?                                !�
���?      �?               @      �?      �?      �?      �?      �?      �?       @                ����'t�?Cw�,��?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?              �?       @���Z��?��d���?      �?              �?              �?      �?       @      �?       @               @       @       @       @       @      �?      �?�}�ɣ��?^͜�ѻ�?                                6���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��*��?�A�m���?              �?                {2~�ԓ�?              �?               @       @                       @       @              �?       @ͤ=����?7�����?      �?              �?      �?3~�ԓ��?      �?       @      �?               @       @               @       @       @      �?        Y7���?�S���J�?      �?      �?      �?        p�z2~��?      �?              �?                       @               @       @              �?       @�yjH��?����~V�?                      �?        Zas �
�?      �?       @      �?                       @       @       @       @      �?      �?        {B���?�	� �?      �?              �?        ?���@��?      �?       @      �?                                                              �?       @�k�.M��?Ѹ��H��?      �?              �?              �?      �?              �?                       @               @       @              �?       @�<݌S�?.F����?                              �?              �?                       @       @               @                              �?       @ٴ��I��?D�z'ys?      �?                      �?��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?��Z#PB�?      �?              �?      �?e�v�'��?      �?       @                       @               @       @              �?      �?       @���S��? �E|��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�? ��?�>      �?              �?      �?�K=��?              �?                                       @       @               @      �?       @�����f�?���U<N�?      �?                        ?���@��?      �?                                                       @                      �?       @�0%fK�?
,�>s��?      �?      �?                p�z2~��?      �?       @                       @               @                       @                ��U�?ʰ�,03�?              �?                �'�K=�?      �?       @      �?               @       @               @       @              �?       @�����?���=�?                                �
��V�?      �?                       @       @                                                       @n��W�?
:��`6�?              �?                ��RO�o�?              �?                                               @       @              �?       @�@ʾ���?�SQ�?      �?              �?        v�'�K�?      �?       @      �?       @               @               @       @       @      �?      �?g�����?�����?      �?                        F���@��?      �?                                                       @                              @؋�ߵN�?}P�7�Ť?                                �]�����?      �?              �?       @                       @               @              �?       @B����?�U\:��?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                        ����[�?:�Z3F�?                      �?      �?��Vؼ?      �?                       @       @       @       @                                      @I!�i��?&���?      �?              �?      �?�@�6�?      �?       @                       @       @               @              �?                      �?�����?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?-h#���?����q�?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?��N�ԑ?����>�?                      �?        (�K=�?      �?       @      �?                       @               @       @      �?      �?       @۴��I��?wv���?      �?              �?        �o�z2~�?      �?                               @       @       @                       @      �?      �?mu����?�_�\H��?      �?                        ���V؜?      �?              �?                                                              �?      @�l	�Y�?��xI�?                      �?        H���@��?              �?                                               @                      �?        Y�՘H�?w�V̓��?              �?      �?        H���@��?      �?              �?               @       @                       @                        Z;��V�?��|_�?      �?              �?              �?      �?       @               @       @       @       @                       @              @S�����?�U۾��?                      �?      �?      �?      �?       @      �?       @                                               @                ����[�?�) �z�?                              �?�ԓ�ۥ�?      �?       @               @                                                              @6A .�?[�>kż?              �?                �K=��?      �?       @                       @                                                       @]!ї�V�?D�ڰ�_�?      �?              �?        �'�K=�?              �?                       @       @       @       @       @       @      �?        ��C���?�����?              �?                	��V��?      �?       @      �?                                       @       @              �?       @���.�?S8� �y�?                      �?        3~�ԓ��?      �?       @      �?               @                                              �?        ��'�?���4��?                                �ԓ�ۥ�?      �?              �?                                                              �?       @ї�V�i�?s}'�;��?              �?      �?        (�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?       @B6w\I`�?��`��j�?      �?                        >�]���?      �?                               @       @       @       @       @       @      �?      �?��Z�<�??@�ਬ�?                                �z2~���?      �?              �?               @                               @              �?       @l	�Y �?��"]v�?      �?              �?      �?���V،?      �?              �?       @                               @       @                       @��vA�?5H0ʉ�?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?              �?      @nC��x�?�7�!\��?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?              �?      @����'t�?�G�O��?      �?      �?                �K=��?      �?       @      �?                                                              �?      @����J�?mϮvD��?                      �?      �??���@��?      �?              �?                                       @                      �?      @��䶺O�?L�T��?      �?              �?      �?P�o�z2�?      �?       @      �?               @                       @       @      �?      �?      �?/��:]�?��e�g��?      �?              �?      �?(�K=�?      �?              �?       @       @       @       @       @               @      �?      �?�ht3Na�?�z�o��?      �?      �?      �?        �
��V�?      �?       @               @       @                                      �?              �?ٴ��I��?Qv��Y�?                                �'�K=�?      �?       @      �?               @                                              �?       @~5&���?�t=O%�?              �?                6��9�?              �?                                                       @              �?       @Sb����?n-��_�?      �?                        ���V؜?              �?                                       @                                       @���J�?zK��F�}?              �?      �?        (�K=�?      �?       @      �?                                                       @      �?      �?�B�]�F�?w:,����?      �?      �?                ��RO�o�?      �?              �?                                       @       @                      �?��ǰ2��?���Nl�?      �?      �?      �?        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?m+�oM�?Y�/C�k�?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @1[�yj�?n� ��k�?                      �?      �?�ԓ�ۥ�?      �?       @      �?       @               @                              �?                #���?O�D%��?      �?              �?      �?�'�K=�?      �?                       @       @               @                      �?              @��U�?F��IZ��?                      �?        �ԓ�ۥ�?              �?                               @               @                      �?       @D�%��}�?ЙǄ;�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?-h#���?ܡ�T��?      �?                      �?                      �?                       @                                              �?      @�r@��?cw�^$�W?                      �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?$�$0�	�?��Ʃ�?      �?                                      �?              �?                                                              �?       @�vAIE�?�!��}�w?      �?                      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                        ����'t�?�0;��?                      �?      �?6���?      �?                                                                      �?      �?      @��j1v�?3H���?      �?              �?        ���Vج?      �?              �?                       @               @       @              �?       @�Gm?C�?X���WQ�?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?w	ܡ�{?      �?              �?        ��ۥ���?      �?       @               @       @       @       @       @       @       @                 J�hY�?2���?      �?                      �?���V؜?      �?                                                       @                      �?      �?E�*�A6�?��fy͑?      �?              �?      �?�o�z2~�?      �?       @      �?                       @               @               @      �?      �?R��'��?�jA���?      �?              �?      �?�K=��?      �?                       @       @       @               @       @       @              �?፿Po�?$�"/���?      �?                        {2~�ԓ�?      �?       @      �?                       @       @       @       @                        Y7���?;�a�Y`�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @M:'>��?b:���9+?      �?      �?                ���.�d�?      �?       @      �?       @       @                       @       @              �?        �mZq�$�?h�D���?                      �?              �?              �?               @       @       @                       @       @      �?       @��̱���?P�u(�N�?                                              �?               @      �?      �?      �?      �?      �?      �?              �?        ]����`�? <���9?      �?              �?        3~�ԓ��?      �?              �?       @       @       @       @       @       @       @      �?      �?$����>�? �^&��?                                              �?              �?                                                              �?       @��w����?˲T dQx?      �?                        ���Vج?      �?       @      �?               @       @                                      �?       @ J�hY�?�i;��?                                P�o�z2�?      �?                       @               @                              �?      �?      �?�ߚ ��?��b�W �?      �?      �?      �?      �?v�'�K�?      �?       @      �?                       @               @       @              �?      �?�۴���?fS��:�?      �?                        3~�ԓ��?      �?       @      �?               @       @               @       @       @      �?        �:Blӊ�?��[4�?      �?              �?        ��ۥ���?      �?              �?               @       @       @       @       @       @      �?       @5&����?4o%��?      �?              �?        p�z2~��?      �?       @               @                       @                      �?      �?       @�n�)L��?r�'�ԝ�?      �?                        P�o�z2�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �^W-��?|���b��?              �?      �?      �?(�K=�?      �?       @      �?               @       @       @       @       @      �?      �?       @� ����?0���,��?      �?              �?      �?��ۥ���?      �?       @      �?       @       @       @       @       @       @       @      �?        ��(��|�?H��_��?                      �?              �?      �?       @      �?       @       @       @       @       @               @      �?        e����I�?�r�����?              �?                ?���@��?      �?       @                                                                              @�I�:Bl�?)�`N��?      �?      �?                e�v�'��?              �?                       @       @               @       @      �?      �?       @#��~���?ܺ�����?      �?                      �?���.�d�?      �?              �?               @               @       @       @              �?      �?9�)1[��?�,ߙ��?              �?      �?        ���Vج?      �?       @      �?               @                                              �?       @�����?�W�+�ؤ?      �?              �?      �?�K=��?      �?       @      �?               @       @               @       @      �?      �?       @��Ͽ�?�
p6a��?              �?                �@�6�?      �?              �?                                       @       @                        +�oM��?�EIg�d�?      �?              �?      �?�K=��?      �?       @      �?               @                               @              �?        �r�9ֳ�?��b�v�?      �?                        �z2~���?      �?                                                       @       @      �?      �?        @�MF��?A�a<��?                      �?        ���.�d�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����'t�?�C�j��?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�፿Po�?��Ur�?                                $Zas �?      �?       @      �?       @                               @                      �?        R��'��?��l�z�?      �?                        F���@��?      �?              �?                                                              �?       @'#��~��?< X��?                              �?Zas �
�?      �?              �?                                       @                      �?       @�����?�G�n�?      �?                        ���V،?      �?                       @               @                                      �?      @xwwwww�?� Co8X�?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @]����`�?�4Znex�?      �?                        �@�6�?      �?              �?                       @                       @                       @y4��0�?�]#ﲹ?      �?                      �?F���@��?      �?                                                                                      @����e�?�:��?      �?      �?      �?        �'�K=�?      �?                                       @       @               @              �?      �? .�c�?<��䠰?      �?                        �
��V�?      �?              �?               @               @       @              �?      �?        �`ph>�?�b�4�?                                ���@��?      �?              �?               @               @       @       @       @      �?      @:'>���?Z����?                      �?        [as �
�?      �?              �?               @                               @              �?        �'�F7��?m��$9��?      �?              �?        F���@��?      �?              �?                                                              �?       @�vAIE�?���y��?                      �?      �?�6��?      �?                       @       @                                                       @,u�ئ�?��/�b�?              �?      �?        3~�ԓ��?      �?       @      �?                       @                                              @���Up�?�(:Q��?      �?              �?      �??���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�%��}�?>;�:�w?      �?              �?        �@�6�?      �?       @                               @               @       @      �?      �?       @�HT�n�?'4�Ջ�?      �?              �?        ��V��?      �?       @               @               @       @               @       @                �.M��o�?W%�*&"�?      �?              �?        �6��?              �?               @       @               @       @       @       @      �?        ٴ��I��?o�C���?      �?              �?      �?��ۥ���?      �?       @      �?               @               @                       @      �?       @y4��0�?a��?                                ���V،?      �?              �?                                       @       @              �?       @���T��?�~�N��?      �?              �?      �?�
��V�?      �?       @      �?                       @               @                      �?      �?���T��?*���x��?      �?              �?      �?���V؜?      �?              �?       @       @                       @                               @t3NaJ��?\��qU!�?                      �?      �?{2~�ԓ�?              �?                       @                       @       @              �?       @���f���?J�_���?                      �?      �?�D+l$�?      �?                                       @       @       @              �?      �?       @F��s�?+eΥ0�?      �?      �?                              �?              �?                                                              �?       @�7�B�]�?���x?      �?              �?              �?      �?       @      �?               @       @       @       @       @       @      �?      �?�n�Wc"�?M=<V���?      �?      �?                ���V؜?      �?       @      �?               @                                              �?       @፿Po�?�����d�?      �?                                      �?              �?                       @               @                      �?       @<��u�4�?p��I�7?                                e�v�'��?      �?              �?       @       @                       @       @      �?      �?      �?��_���?3A2���?      �?                        �@�6�?      �?                       @               @       @       @       @                      �?���Y;�?P��~q�?                                                      �?               @                                                              @�\d����?^��HY�T?      �?      �?      �?        �z2~���?      �?              �?                                               @              �?       @*L����?�%4���?                                              �?                       @                                                      �?      �?K���S�?'�d��+l?                                ��RO�o�?      �?              �?               @       @               @       @      �?      �?      @��'t �?��e
�"�?      �?                        �@�6�?      �?       @      �?               @       @               @       @              �?       @�oM���?h��l���?      �?      �?      �?              �?      �?       @      �?       @       @       @               @       @       @      �?        �C��?��=��-�?      �?                        ���Vج?              �?               @       @       @       @                              �?      @_ph>��?d
����?      �?              �?        e�v�'��?      �?       @      �?               @       @               @       @              �?       @��0%f�?C揮k�?                      �?      �?�K=��?      �?       @                               @       @               @       @      �?        X-�r�?�t*����?      �?                        !�
���?      �?       @               @                       @                      �?              �?Ήo���?�=�V�?      �?                              �?      �?       @      �?               @       @               @       @       @      �?       @��8�)1�?G�Zln�?      �?                        H���@��?      �?       @      �?               @       @               @       @              �?        ��-�<5�?�\�k��?      �?      �?                �ԓ�ۥ�?      �?       @      �?                                       @       @              �?       @��f��?�@�����?      �?      �?      �?        ��V��?              �?                       @       @       @       @                      �?       @��e0
8�?�$i@��?      �?                      �?�'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @�r@��?@?��_
�?      �?      �?      �?        3~�ԓ��?      �?       @      �?               @       @                       @              �?       @����?��_��?                                �V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?       @$�$0�	�?�epؓ �?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�፿Po�?L���ξ?              �?                                      �?                                               @                      �?       @�5A .�?�PC_B�`?                      �?      �?P�o�z2�?      �?       @      �?               @       @                               @      �?      �?a�:�?�9>��&�?                      �?      �?ܥ���.�?      �?                       @               @       @       @              �?                K��a�?��Ǉ�0�?                      �?      �?Zas �
�?      �?                       @       @               @               @       @                _ph>��?Ky&Hf0�?                                ��Vؼ?      �?              �?                                       @       @              �?        �?y4��?���]�?      �?                        �'�K=�?      �?              �?                       @               @                               @ J�hY�?ePm��?                      �?        �o�z2~�?      �?       @               @       @               @       @       @       @      �?       @Ô�-�<�?�6���?      �?              �?        ���.�d�?      �?              �?               @       @       @       @       @      �?      �?      �?��E�X��?�^I_��?                      �?      �?�o�z2~�?      �?       @      �?               @               @       @       @      �?      �?      �?g�����?�*����?      �?                         �
���?              �?               @                       @       @       @      �?              �?�
n���?���#��?                                e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @              @Y�)L�ْ?�#8�U�?      �?                        ���V؜?      �?       @      �?                                                              �?       @�u�b���??��o �?      �?                      �?�'�K=�?      �?                                       @       @                      �?              �?��J�ć�?dB�b���?      �?                        !�
���?              �?               @                       @               @              �?      �?�r@��?u�����?      �?                        ��RO�o�?      �?                       @               @       @       @              �?              �?�vAIE�?킸ar0�?      �?                                      �?              �?                                               @              �?       @�I�:Bl�?^\�Wa�|?      �?              �?      �?�6��?      �?       @      �?               @       @               @                      �?       @�<݌S�?���[���?                                H���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?����[�?7r[��S�?                                �o�z2~�?      �?                       @                       @               @       @      �?      @UH�%���?���!&E�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�d�Q�ϐ?��<��?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        Y�)L�ْ?��9�z��?      �?              �?      �?v�'�K�?      �?              �?       @       @       @               @       @      �?      �?        3��g�?n}�����?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?E�(Ţe�?vG���Q?      �?                      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @                ,1[�yj�?pQݖ?      �?              �?        �]�����?      �?              �?       @       @       @                                      �?      �?J̖p���?zw�;�?                                ?���@��?      �?       @                                       @       @                      �?      @ .�c�?"���{��?      �?      �?      �?        �RO�o��?      �?              �?               @       @               @       @      �?      �?       @�6��`�?�2�R��?              �?      �?        ��V��?      �?       @      �?       @       @       @               @       @              �?      �?x�/���?��ҩ\��?                      �?      �?$Zas �?      �?       @      �?               @       @               @       @              �?        [�KS}��?��-&�f�?                      �?      �?���.�d�?      �?       @      �?               @       @                       @      �?      �?       @/������?��#��?                      �?      �?���.�d�?      �?               @      �?      �?      �?      �?      �?      �?      �?                -h#���?Q'a�w�?      �?              �?        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?n��W�?t�����?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?              �?       @Z��2�?L�9�(�0?                                	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?                �d�Q�ϐ?R9+�?��?      �?      �?      �?              �?              �?               @       @       @       @       @       @       @      �?      �?Ň7�B��?���?                                �@�6�?      �?       @      �?       @                                                      �?       @����[�?j��g��?                      �?        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?                ś�8j��?�M{��?      �?                        �'�K=�?              �?                                                              �?      �?      @�d�Q�ϰ?k` �e��?      �?                                      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @)g��1�?徢�qG?                              �?��V��?              �?                       @               @       @               @              @)g��1�?}"�$g��?      �?      �?      �?        �D+l$�?      �?       @      �?                               @       @       @              �?       @���?A��h�?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @!�iŽ�?��`Y��?      �?              �?        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?       @F��1��?��#��?                              �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?Y�)L�ْ?�kѥ�{�?      �?                        ,l$Za�?      �?              �?                                                                      �?U�����?�n���?                      �?        p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?���C�?`����i�?      �?                        ��.�d��?      �?       @      �?       @               @       @       @       @       @      �?       @�MF���?��$�?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?E�(Ţe�?Go�L�?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @       @                 �&#���?� ����?      �?              �?        Zas �
�?      �?                       @       @               @       @       @       @      �?      @O�)���?_uS�2v�?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?�9�(� ?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�L�5A �?�?Y�/?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?               @       @       @       @       @       @      �?       @ۙ�ǰ2�?z�S��?                                ��V��?      �?       @      �?       @                                       @              �?       @�ߚ ��?0��|���?      �?              �?      �?��Vؼ?              �?                       @                                              �?       @˲
n�ͽ?9^��1�?                      �?        �@�6�?      �?                       @               @       @       @       @      �?              @m$���?x<��?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�����`�?���jj�?                      �?        �ԓ�ۥ�?      �?              �?       @       @               @       @       @      �?      �?      �?�]�FR�?Bǁy��?                      �?      �?      �?      �?                       @       @       @       @               @       @      �?       @,�����?7z�')E�?                      �?      �?�@�6�?      �?       @               @       @       @               @              �?      �?      �?&`��"�?=�]ݒ��?      �?              �?        �
��V�?      �?       @      �?       @       @                       @                      �?       @��C���?Ś'�F�?                      �?        ܥ���.�?              �?               @               @                       @              �?        �����9�?����g�?              �?      �?        �K=��?      �?       @      �?               @       @                       @              �?       @��s��2�?UZC<���?      �?      �?      �?                      �?       @      �?                                                                       @j�����??ښo;z?                                �@�6�?      �?              �?               @               @       @       @       @      �?        ��w�ӥ�?l�]6��?                                �6��?      �?       @                       @               @               @                      �?S�����?��s�yz�?                      �?      �?��V��?      �?       @      �?               @       @       @       @       @       @      �?      �?����w�?߿R�ͯ�?                      �?      �?      �?      �?       @               @       @       @       @       @       @       @                #��~���?�U�����?                                Zas �
�?      �?       @               @       @       @       @       @       @       @               @h{����?%s����?      �?                        [as �
�?      �?       @                       @               @       @                      �?       @�d�Q���?ysT�&��?                                ܥ���.�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                I`�:�?�IbBN��?              �?                �ԓ�ۥ�?      �?              �?               @                                              �?       @�6��`��?��Z���?                      �?      �?�z2~���?      �?                               @               @                      �?      �?      �?^!ї��?T#aI��?      �?                        ��Vؼ?      �?              �?                                                                      @���"X~�?��_h޲?              �?      �?        �RO�o��?      �?       @      �?       @       @       @       @       @       @       @      �?        �:]��#�?�IbBN��?      �?              �?      �?�ԓ�ۥ�?      �?                       @       @               @       @       @       @                7w\I`��?��|��e�?                                �]�����?      �?       @      �?               @       @               @       @       @      �?       @M�cX�~�?G��(���?      �?              �?      �?��ۥ���?      �?                       @       @       @       @       @       @       @                b�(Ţe�?���SP2�?                                              �?              �?       @                                                              @���H*�?sn:Oo�z?                              �?�]�����?      �?              �?       @       @               @       @       @      �?      �?      �?�*g���?��[����?      �?              �?        P�o�z2�?              �?               @               @               @       @       @      �?        ��7q��?9qR_]��?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @�d�Q�ϐ?��nh:�?      �?              �?      �?6��9�?      �?       @               @               @       @                       @      �?      �?8j��^�?�q`^���?      �?                        ܥ���.�?      �?       @      �?               @       @               @       @      �?      �?      �?)����?�MP��?                      �?      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?       @              @�]�FR�?B���Rbo?                                e�v�'��?      �?       @      �?               @       @               @              �?      �?        &���[�?������?                      �?      �?[as �
�?      �?       @                       @               @       @       @       @                ��r�9��?�F��G�?                      �?      �?�D+l$�?      �?       @      �?                       @               @       @              �?       @��_���?'�1m�[�?                      �?      �?��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?!�iŽ�?��KA*�?                      �?        ���V،?      �?       @      �?                       @       @       @       @              �?       @A���Kn�?�V
u�w�?                      �?        P�o�z2�?      �?       @               @       @       @       @       @       @       @      �?       @����c�?=����?                                ��V��?      �?              �?               @               @                      �?      �?        �`�AQ��?���s��?      �?                        ��V��?      �?       @      �?       @                       @               @      �?               @������?����W�?                      �?      �?v�'�K�?      �?                       @                               @               @      �?       @<�RG�m�?�yz��`�?                      �?        �@�6�?      �?       @      �?       @                       @       @                      �?      �?Aʾ����?=�h���?                      �?      �?3~�ԓ��?      �?                       @       @       @       @       @               @              �?x�ӥ�>�?�=G�P�?      �?              �?      �?�
��V�?      �?              �?               @               @                                       @)�tN|x�?㥉�)�?                                �K=��?      �?                       @       @                                      �?              @jL�*g�?w�!���?                      �?      �?(�K=�?      �?       @               @       @       @       @       @               @                �j1v��?ӡ��c#�?      �?              �?        ���V؜?              �?                                                                              @)g��1�?�,V�a|?      �?              �?        3~�ԓ��?      �?       @                       @               @               @       @              @�e0
84�?�/k�!�?              �?                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?��%xH+�?      �?                        ���V؜?              �?                               @               @                      �?      @Z�KS}��?��t�?                      �?      �?6���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�'�F7�?Lp����?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @      �?      �?xwwwww�?ߖ �P[�?      �?              �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����'t�?~�杭��?              �?      �?              �?      �?       @      �?       @               @       @       @       @       @      �?      @�n�Wc"�?�����?      �?              �?        (�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                b��1��?��K0�?                      �?      �?      �?              �?               @               @               @       @       @      �?      �?�G�Ɉ��?��{q��?                                �'�K=�?      �?       @                                                                      �?       @�`�AQ��?���߄�?              �?                SO�o�z�?      �?       @      �?                                       @                      �?       @0��m$�?������?      �?                      �?              �?       @      �?                                       @       @              �?       @�H*���?����4��?      �?              �?              �?      �?       @               @       @       @       @               @       @      �?        ]��#�d�?o鵽��?      �?              �?      �?��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?���5��?                      �?      �?�ԓ�ۥ�?      �?       @               @       @               @       @              �?              �?E_r[ݧ�?�N����?      �?              �?        SO�o�z�?              �?               @                               @                      �?        Z�KS}��?��)[��?              �?                ���.�d�?      �?                       @       @               @       @               @      �?      �?��6���?"z�?              �?                      �?      �?       @      �?               @       @       @       @       @       @               @Ň7�B��?��3C�?                                 �
���?              �?                               @               @       @              �?      �?���7q�?�\��i��?      �?      �?                              �?              �?                                       @                      �?       @��&`�?���:�|?      �?              �?      �?�V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?F��1��?��˻��?      �?              �?      �??���@��?      �?       @      �?               @       @                                      �?        y4��0�?[YU)�ܤ?                                �o�z2~�?      �?       @      �?       @       @       @                              �?      �?       @�a/��?q�4/�?      �?              �?      �?F���@��?      �?                                                                                       @ꏗ�(��?Sw���?                      �?        ��RO�o�?      �?              �?                       @               @       @      �?      �?        �g�L�c�?:<�M�d�?                      �?        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?�R��e?      �?              �?        ��.�d��?      �?       @               @       @       @       @               @      �?      �?      �?�X����?��;K��?                              �?              �?              �?                                               @                       @���Y;�? �|��I|?      �?                        F���@��?      �?              �?       @                                                      �?      �?*g���?��Hl��?      �?              �?      �?6���?      �?       @      �?                                       @               @                jŽ�,u�?�ߟf3��?                      �?      �?      �?      �?       @      �?       @               @       @       @       @       @              @�����f�?�S{[���?      �?              �?        �]�����?      �?              �?       @               @       @                      �?      �?        ~5&��?������?      �?                        p�z2~��?      �?       @      �?               @                       @       @              �?        �p����?V��/��?      �?                        ���V؜?      �?              �?                                       @                               @�I�:Bl�?�^� f�?                                �z2~���?      �?       @               @                                                               @ J�hY�?s�=�,�?              �?      �?      �??���@��?      �?                                                                                       @*g���?�J-�<�?      �?              �?      �?!�
���?              �?               @       @       @               @       @      �?               @���+$�?�jj���?      �?                        ��ۥ���?      �?       @      �?                       @       @                       @      �?      �?݌S���?���2���?      �?      �?      �?        ��V��?      �?       @      �?       @       @                       @               @      �?      �?�X�ڙ��?%�x-��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @F��1��?��ֺ�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      �?�U�����?��8�g��?                                              �?                                                       @                      �?       @�5A .�?�7x��p?                      �?        ���Vج?      �?              �?       @               @                       @              �?      @�&#��~�?E?����?      �?                        F���@��?      �?              �?               @       @                                      �?       @A .��?��:�x3�?              �?                ��RO�o�?      �?       @      �?               @       @               @       @              �?       @�+$���?��"�vW�?                                Zas �
�?      �?              �?               @                                                        ��8j��?
�`���?      �?              �?        �V�H�?      �?       @      �?               @       @               @              �?      �?       @�<݌S�?��<����?                                !�
���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        m+�oM�?�/(W0�?      �?                      �?�D+l$�?              �?                                               @       @              �?       @K�*g��?�o��	�?      �?              �?        �o�z2~�?      �?       @      �?                       @       @       @       @       @      �?        `��"s�?o^���t�?      �?                        �@�6�?              �?                       @               @                              �?       @��D)�?�Ԙ:�?      �?              �?      �?{2~�ԓ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��N�Ա?� T[o0�?                                �ԓ�ۥ�?      �?              �?                       @       @       @       @      �?      �?       @����?]����?                      �?        ���@��?      �?       @      �?       @       @               @       @       @              �?        H���<�?3H�Y��?                      �?      �?�
��V�?      �?       @               @               @       @       @       @       @      �?        �vAI�?��g!�?              �?      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?Dz�rv�?��>[�?      �?                        ���V،?      �?       @                       @                                              �?      @ J�hY�?�2�R���?      �?                        6��9�?      �?                                       @       @                              �?      �?jL�*g�?�9�[�?                      �?      �?              �?                                       @                                              @�%��f��?�|�:�m?                                ���V؜?      �?              �?                                                              �?       @��w����?�UO��?                      �?      �?���Vج?      �?              �?               @                               @              �?       @.2�z���?ɱ��Ŧ?                      �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @              @F��1��?,Uwm�y�?                      �?      �?>�]���?      �?       @               @                               @              �?                dsǕ��?M�F���?                      �?        e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?n��W�?R��R�?      �?                        e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @              @��N�ԑ?O\���?      �?              �?        ��ۥ���?      �?       @               @       @       @       @               @       @              �?g��}���?���?      �?                        6��9�?      �?       @                                               @       @                      @�l	�Y�?0�LR�?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�'�F7�?m>sR�?                                �z2~���?      �?              �?       @                                                      �?        �N���?�@�Z���?                                ���V،?      �?              �?       @       @                       @                      �?       @F�*�A6�?����a��?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�X����?K�b�Zs?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?                      @]����`�? <���9?      �?              �?        	��V��?      �?              �?                       @               @       @      �?      �?        �Y;���?�g�m.�?      �?              �?              �?      �?       @               @       @       @       @       @       @       @      �?      �?��O�n�?�<�L?3�?      �?              �?        ���V؜?      �?                                       @       @                              �?      @ͤ=����?�C��e
�?      �?                        ���Vج?      �?       @      �?               @       @               @       @                       @���_���?��y�ek�?      �?      �?                �o�z2~�?      �?       @      �?               @       @       @       @       @      �?      �?        F��s�?-|����?      �?                      �?�'�K=�?      �?       @      �?               @       @       @               @      �?              �?���?y4�?�E����?                                              �?                               @                                              �?       @K���S�?'�d��+l?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?      �?              @�0[�yjv?              �?                        ���V،?      �?              �?                                                              �?      �?ї�V�i�?���c�?                                F���@��?      �?       @      �?                                               @              �?       @l	�Y �?���1�?                                6��9�?              �?                       @               @                                       @���@���?�HY��?      �?      �?                �'�K=�?      �?       @                       @       @               @       @       @      �?        ~5&���?�����Q�?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @8�]�FR�? ���WYw?      �?              �?      �?v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?��N�ԑ?+
��?      �?              �?        [as �
�?      �?       @                               @       @       @       @      �?      �?      @���Up�?d��k�4�?      �?                        [as �
�?      �?                                       @       @                              �?       @
84���?W�"'�?      �?              �?      �?	��V��?              �?               @               @               @              �?              �?�r@��?YRgض?      �?              �?        !�
���?      �?       @      �?               @       @               @       @      �?      �?        ճv&�1�?��UZC<�?      �?                        ��RO�o�?      �?              �?               @               @                              �?      @r�g�L��?xp�7��?                      �?        $Zas �?      �?              �?                       @       @                              �?      @�����?ON��W��?                                6���?      �?                       @       @       @       @                       @      �?      �?@�MF��?���*)��?      �?              �?        H���@��?      �?              �?                               @       @       @              �?      �?��.h#��?:Z~[!�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @-h#���?��??              �?      �?        6��9�?      �?              �?                       @       @       @                               @��,u���?�R��?      �?              �?      �?�ԓ�ۥ�?      �?                       @       @       @                               @      �?        <�RG�m�?6V��	��?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?��;�l|~?      �?      �?      �?                      �?       @      �?                                       @                      �?       @�����?xjD",�?      �?                      �?��ۥ���?      �?                       @       @       @       @       @               @      �?      �?�X���?*��R�?                                �'�K=�?      �?       @      �?       @       @       @               @       @       @      �?        �U:'�?��ㅝ��?                                Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?,1[�yj�?c���Y�?      �?      �?      �?        ,l$Za�?      �?       @      �?                       @               @                      �?       @��ߵN��?y��	��?                                H���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?Q6��$�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @���@��?�ppTV�)?                                ���V،?      �?              �?                                               @                       @�F���?xv6���?      �?              �?      �?	��V��?      �?       @      �?                                       @       @              �?       @����_��?z�A���?                      �?      �?6���?      �?       @               @               @       @       @               @              @G��q
S�?��s<�?                      �?        Zas �
�?      �?       @      �?               @               @               @       @      �?        |]�;�?XYHK��?                      �?        6��9�?      �?       @      �?                       @                                      �?      �?L���S�?�i3a��?              �?                6��9�?      �?       @      �?                                                              �?       @#�6��w�?�D�����?                                F���@��?      �?       @      �?                                                              �?       @k� 6\.�?f����?                                �ԓ�ۥ�?      �?       @      �?               @               @                                      �? J�hY�?�i�kMh�?                      �?      �?�ԓ�ۥ�?      �?       @      �?       @       @       @       @       @              �?      �?      �?����Z��?�h�XO��?                      �?        �@�6�?      �?       @      �?               @       @               @       @              �?       @���_���?��\��?      �?      �?                $Zas �?      �?       @      �?               @                               @                       @j��|��?�w�!��?                                �'�K=�?      �?              �?       @       @                       @       @              �?      �?u�4�G��?��F�o��?      �?      �?                �z2~���?      �?       @      �?                       @               @       @              �?       @�E�X���?�����r�?      �?                        �'�K=�?      �?       @      �?       @                               @       @              �?       @�;�$0��?��dO!��?                      �?      �?��V��?      �?       @               @       @       @       @       @       @       @      �?      @��ǰ2��?D�J~@��?                      �?      �?��ۥ���?      �?                       @               @       @       @       @       @      �?      �?��-�jL�?)j�K��?      �?                        ���V؜?      �?       @      �?                       @               @       @              �?        ωo���?8G'��?      �?              �?      �?P�o�z2�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�rv��?��kh���?      �?      �?                ��V��?      �?       @      �?               @       @                                      �?      �?�'�F7��?&�����?      �?                        F���@��?      �?                                       @       @       @                                ��Z�KS�?m���<�?      �?                        �ԓ�ۥ�?      �?              �?               @       @               @       @      �?      �?        �5\.2��?A[�����?                      �?      �?��.�d��?      �?       @      �?       @       @       @                       @                        ��	�p�? "��^�?                      �?      �?�V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @8�]�FR�?�G��Ժ?      �?              �?        �z2~���?      �?       @      �?               @       @               @       @              �?        Q���\�?G����?      �?                        F���@��?              �?                                                              �?      �?      �?��*��?��N��4�?                                              �?              �?                       @                                               @���H*�?sn:Oo�z?                                              �?              �?                                                              �?       @>�/�Q�?U�9��w?      �?              �?      �?P�o�z2�?      �?                       @       @       @       @                       @              �?��>�MF�?����?                      �?      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?O�)���?�+� n�?      �?              �?      �?�RO�o��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �X����?�x�q"}�?      �?              �?      �?F���@��?      �?                                       @                                               @Y���d�?�Ѹ����?                      �?      �?e�v�'��?      �?       @                       @       @                               @      �?        �^<��u�?Gɶ�7��?      �?              �?        (�K=�?      �?                       @       @               @               @       @              @;��V��?����C'�?      �?              �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ����'t�?�h�v,-�?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?G�S�y_�?                      �?      �?��ۥ���?      �?       @      �?               @       @               @                      �?        ��B�/�?=����e�?      �?              �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @���f�´?z�H�9�?      �?                        �
��V�?      �?       @      �?                                       @       @              �?       @fK8O��?u&*q�?                                �@�6�?      �?              �?       @                                                               @m$���?r� Co8�?              �?                �]�����?      �?              �?       @       @                                                       @8q��3�?���) ��?      �?              �?      �?��.�d��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?9�%��}�?��\��?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�X����?���:�t?                      �?      �?>�]���?      �?       @      �?                       @               @       @      �?      �?      �?!ї�V��?}jL� L�?                                �o�z2~�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?���Y;�?r]����?                                ���Vج?      �?       @      �?                       @               @       @              �?       @����e0�?�A�A�?      �?      �?      �?        ��V��?      �?       @      �?               @       @               @       @      �?      �?        3��g�?Ԫ'�?      �?                        ��RO�o�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?�r@��?`�y�Q�?      �?              �?        SO�o�z�?      �?       @      �?               @       @       @               @              �?       @�E�X���?%��k�?      �?              �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        �X����?�1?��$�?      �?      �?                $Zas �?      �?       @      �?                                       @                      �?       @����?))EC��?      �?      �?                �'�K=�?      �?              �?                                                              �?       @K��a�?~���]�?      �?                      �?�ԓ�ۥ�?      �?       @               @       @       @       @       @               @      �?      �?�ti��|�?���?�?      �?              �?        ��.�d��?      �?              �?       @                               @                               @�W���?Dj��?      �?              �?        ���.�d�?      �?              �?       @                                                      �?      @���G���?���r���?      �?                        �K=��?              �?               @                       @       @               @               @���U�?{d��?      �?                        e�v�'��?      �?                       @       @               @       @                      �?      @X-�r�?�)@��?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                        �X����?�ؐ^�?      �?              �?      �?6���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @�%��}�?�I���?                                ��Vؼ?      �?       @      �?                                               @              �?       @�q
Sb��?x��,�?                                ���Vج?      �?       @      �?                                                                       @x�ӥ�>�?�O��T�?      �?                        �ԓ�ۥ�?      �?       @      �?                                       @                                �H*���?���
p�?      �?              �?      �??���@��?      �?       @                                                                      �?       @jg����?ľl�o�?      �?              �?      �?F���@��?      �?       @                       @       @       @       @                      �?       @�<�^�?��,C�?              �?      �?        �]�����?              �?                       @       @               @       @                      �?.������?x�3�(�?      �?                        ���Vج?      �?              �?                                               @                      @?^��C�?p�"�?                                �RO�o��?      �?              �?       @               @       @       @       @              �?        �e� ��?on�����?      �?      �?      �?        �D+l$�?      �?                               @                                              �?        +���?y�?��&��H�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�X����?,g��	�?                      �?        (�K=�?      �?       @      �?                       @               @       @      �?      �?       @[�yjH�?��$T϶�?      �?              �?      �?���@��?      �?                                                                      �?      �?        q%�yO��?�t`�V�?      �?              �?        �V�H�?              �?               @               @       @                       @              �?�~k� 6�?*9�\���?      �?              �?        Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                n��W�?1+�^�r�?                      �?      �?�
��V�?      �?              �?                                                       @      �?      �?b����,�?$��M=�?      �?              �?      �?      �?              �?               @       @       @       @                       @              �?)g��1�?�"���?      �?      �?      �?        �D+l$�?      �?              �?       @       @       @                              �?      �?      �?F�X�ڙ�?�Ntm1	�?                      �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              @m+�oM�?_I���?              �?                F���@��?      �?                       @                                                      �?       @݌S��?\��e��?      �?              �?      �?��V��?      �?       @      �?                       @       @       @       @       @      �?        �����U�?��ϫ�?                      �?      �?���Vج?      �?              �?                                       @                      �?       @B�/����?eb%��?      �?                        p�z2~��?      �?       @      �?               @                       @                      �?      �? J�hY�?�'�ܷ�?      �?                        �K=��?      �?       @      �?       @       @       @       @       @       @      �?      �?        �Y e��?>�����?      �?              �?      �?�o�z2~�?      �?              �?       @       @       @       @       @       @       @              @kH����?�����"�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      �?^��Z��?@9N�O,�?      �?                        p�z2~��?      �?       @      �?               @       @                                      �?        <��u�4�?a��B���?      �?                                      �?              �?                                                              �?      @D)-��?]v�{x?                                p�z2~��?      �?       @      �?               @       @               @       @              �?       @����>�?<��s��?                                ���V،?      �?              �?                                                                       @� �;�$�?E�v�jۇ?                                 �
���?      �?       @      �?                       @               @       @              �?        ����e0�?�+����?                              �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�U�����?�Ҧ����?      �?                        3~�ԓ��?      �?       @      �?               @                                              �?        ���!���?�u���?      �?                        3~�ԓ��?      �?       @      �?       @                       @                                        �Y;���?�S���J�?      �?                        �z2~���?      �?              �?                       @               @       @      �?               @��.h#��?�R���5�?                                              �?               @      �?      �?      �?      �?      �?      �?                      �?�፿Po�?@}m[&?                      �?      �?      �?      �?       @      �?       @       @       @               @       @       @              �?
���O�?�2H���?      �?                                      �?                                                                                      @�}��j�?p~#ĉUi?                      �?      �?F���@��?              �?                                                                      �?       @�bѲ
n�?��Ȏ?      �?                        !�
���?      �?               @      �?      �?      �?      �?      �?      �?       @              @1[�yj�? �Z��>�?              �?      �?        �
��V�?      �?       @      �?                               @       @       @              �?      �?��G��q�?�(ִ8��?                      �?      �?�'�K=�?      �?                                                                                       @+�����?���U�?      �?      �?      �?        $Zas �?      �?              �?               @                                              �?       @��}�ɣ�?zofC�V�?      �?      �?      �?        ���V،?      �?              �?                       @                                      �?       @�J���?���{���?              �?                �@�6�?      �?       @      �?               @                       @       @              �?       @�C��x�?O��R�?      �?                        ,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?���C�?�� �1�?      �?      �?      �?      �?3~�ԓ��?      �?              �?               @                       @       @              �?      @�%��}�?�,�zU��?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?                      @����'t�?�G�O��?      �?              �?      �?v�'�K�?      �?                       @       @       @       @                       @              @3���O�?�#-^�?                      �?        �
��V�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @<݌S��?��VJM�?      �?                                      �?                                                                              �?       @Z��r�?0-V�ai?      �?              �?      �?�z2~���?      �?       @      �?               @       @                       @              �?        q��3���?��@uc�?      �?                         �
���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        �X����?>��PĪ?      �?                        {2~�ԓ�?              �?               @       @       @               @       @      �?              �?Z�KS}��?�P~~�h�?      �?      �?      �?        ���.�d�?      �?              �?       @               @                              �?              �?������?�b`Czu�?                                �K=��?      �?               @      �?      �?      �?      �?      �?      �?      �?               @�፿Po�?Gqm����?                      �?        ��ۥ���?              �?               @       @       @       @       @       @      �?                )$�����?����>�?      �?      �?      �?        ��ۥ���?      �?              �?               @       @       @               @       @      �?      �?��[�՘�?��C���?                                ���V،?      �?              �?       @       @               @                              �?       @�,u�ئ�?��_*>�?      �?      �?      �?        �o�z2~�?      �?       @      �?               @       @               @       @      �?      �?       @Wc"=P9�?ŗTin��?              �?      �?      �?�
��V�?              �?                       @                               @      �?      �?       @R�&#��?�<���ֿ?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?}m[&r?                                �]�����?      �?       @      �?                                       @                      �?        ��Kn���?�����?                      �?      �?�D+l$�?      �?       @                               @       @       @               @      �?        ���q%�?J��D��?                      �?      �?      �?      �?       @               @       @               @                       @              �?��۴��?���(��?                      �?        �'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @��Po��?���Υ?      �?              �?        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        1[�yj�?\�$ȶ?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?       @              @E�(Ţe�?J���q'?      �?                        ?���@��?      �?              �?                       @                                      �?       @Q�E�*��?�K�����?      �?              �?      �?v�'�K�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?��+$��?��X��?                                              �?                                                                              �?      @�'t J�??�{#%i?      �?              �?      �?3~�ԓ��?              �?                       @       @       @                       @                ��V���?�:'���?      �?                                      �?                                                                                       @�����9�?���W�i?                      �?      �?�K=��?      �?       @      �?               @               @       @               @              �?=���&�?mRI4�?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�����`�?��n�X�%?                      �?      �?�@�6�?      �?       @      �?               @       @       @       @       @      �?      �?        �"s�g��?;�ީ�`�?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                �d�Q�ϐ?j�`F<3�?      �?              �?      �?���@��?              �?               @                               @                      �?      �?�L�5A �?;4����?      �?                        ���V؜?      �?              �?               @                               @                       @�H*���?0�����?                              �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?q������?                                              �?               @      �?      �?      �?      �?      �?      �?                       @����'tx? �<$3�>                      �?        �@�6�?      �?                                                                                      @Z��r�?������?      �?              �?        �'�K=�?      �?              �?       @                                                      �?      @�N���?P-#���?      �?              �?      �?F���@��?      �?                       @               @       @               @              �?      �?q%�yO��?t޶L\�?              �?                ���Vج?      �?              �?                                               @                       @L���S�?����>�?      �?                        ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?      �?                8�]�FR�?�E I�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      �?�U�����?r��1֑?      �?              �?      �?���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�?���Z�?                                Zas �
�?              �?               @       @       @       @                      �?              �?�Kn��4�?�Y䣒��?      �?              �?      �?��.�d��?      �?       @      �?               @               @               @              �?        HT�n��?(Tn'��?      �?              �?        ���@��?      �?       @      �?       @               @               @       @      �?      �?       @e����I�?��`�d?�?      �?                      �?�z2~���?              �?               @               @       @                       @              @K|x�/��?�a�ȸ?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @-h#���?�M����?      �?              �?      �? �
���?      �?       @      �?                                       @                      �?       @x�����?�<wuKN�?      �?                        ��RO�o�?      �?                       @                       @                                      @*1[�yj�?F���N�?      �?              �?        (�K=�?      �?       @      �?               @       @               @              �?      �?        ���`p�?p�7�O�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�%��}�?����?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?              �?       @�፿Po�?�!�0�?      �?                        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @                ���@��?���)���?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?[�<��?�<�L?3�?      �?              �?        v�'�K�?      �?       @      �?               @       @               @       @              �?      �?e0
84��?z{PE�?                                              �?                               @                                                       @�Po���?&��=mn?                      �?              �?      �?       @      �?       @       @       @               @       @       @      �?       @�C��?�y�̹�?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @      �?      �?���l	�?_��F���?                      �?        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                       @����[�?���B(�?                                              �?                                                                              �?        ~PT���?B֜�#�h?                      �?        �@�6�?      �?       @      �?       @               @               @       @              �?        A���Kn�?�w"�C�?      �?              �?      �?F���@��?      �?              �?                       @               @       @              �?      @�Y;���?1������?      �?                        �@�6�?      �?       @      �?               @                                              �?       @ e��h�?\�x��?                      �?      �?�K=��?      �?                       @       @       @                              �?      �?      @>|]��?hl�RW��?      �?              �?        �'�K=�?      �?       @      �?                       @               @       @              �?       @�ht3Na�?�Q�I��?                                �'�K=�?      �?       @      �?                       @               @       @              �?       @�p����?vs�e̮�?                                �@�6�?      �?       @      �?                                                                       @��~5&�?0#=�-��?                                              �?              �?                       @               @                      �?       @b�(Ţe�?;�
���?      �?      �?      �?              �?      �?              �?       @       @               @                       @      �?      �?y4��0�?�����?                      �?      �?�
��V�?      �?       @               @       @               @               @      �?      �?        �ئ�N�?$l@4zZ�?      �?                        �ԓ�ۥ�?      �?       @               @       @       @       @               @       @      �?      �?+�d�#�?Ґ �o�?                      �?        �]�����?      �?       @      �?       @       @                               @              �?       @=���&�?n�� �1�?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?               @                       @                      �?       @��7q��?�ؐ^��?                      �?        6���?      �?       @      �?               @       @                       @      �?      �?       @J�hY7�?ۓ�˅��?                                ?���@��?      �?              �?               @       @       @       @       @      �?      �?       @O|x�/��?�����?      �?              �?      �?�o�z2~�?      �?       @      �?       @       @                       @              �?      �?      �?3��l�?Z��HQ�?      �?                        6���?      �?       @      �?                               @                                        7w\I`��?�Qt���?      �?                        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?�X����?C�7�^�?      �?              �?              �?      �?       @               @       @       @       @       @       @       @      �?      �?:Blӊ{�?�DPk��?      �?      �?      �?        >�]���?      �?                       @       @       @       @       @       @       @      �?        o��4�u�?T+�5̾�?                      �?        {2~�ԓ�?      �?       @                       @                                                      �?2��l�?SB3Nfn�?                                ��RO�o�?      �?                               @               @                              �?      @z����"�?��EIg��?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�U�����?;b/��b?      �?              �?      �?�]�����?              �?                       @                                                      �?�S��%�?0���N��?                      �?      �?���@��?      �?       @               @       @       @       @               @      �?      �?        ���w��?�n���?      �?                      �?      �?              �?               @       @       @       @       @       @       @              �?]�FR,�?�b�g.�?      �?                        ���Vج?              �?                                                                              @�c=kgҮ?ƶJ-�<�?      �?                        	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        �U�����?�˨�?      �?                        $Zas �?      �?                                               @                                      @��e0
8�?����Q�?      �?      �?      �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?-h#���?:�\��:�?                      �?        �
��V�?      �?       @               @       @               @                      �?      �?      �?MaJ̖p�?#�~N�m�?      �?              �?        6��9�?      �?       @               @                                                      �?      @�፿Po�?Qu����?      �?              �?        ��ۥ���?      �?       @      �?       @       @       @       @       @       @       @      �?        �R��'�?��]8��?      �?      �?      �?        {2~�ԓ�?      �?                                                               @      �?               @ͤ=����?`H3�G��?      �?                        �z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�?y�S�?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      �?1[�yj�?M3�z�n�?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?�Y;���?�0g�~?                                              �?                                                               @              �?       @����_��?.[�ɎLq?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?E��a�?2�"ml(�?      �?                        �'�K=�?      �?       @      �?               @               @               @                       @��.h#��?�)�-�'�?                                F���@��?              �?                       @                               @              �?      �?K|x�/��?�U$��7�?                      �?      �?Zas �
�?              �?                       @       @       @       @               @              �?$���?���W��?              �?      �?      �?{2~�ԓ�?      �?       @      �?                                       @       @              �?      �?�0%fK�?A�&���?      �?                        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                zyO�0@�?�fQ0��?      �?                        �@�6�?      �?              �?                                                                       @��6���?�xP��?      �?                        ���V؜?      �?              �?               @       @       @       @       @              �?       @_�ti���?ۄ��n��?      �?              �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @h#���?l
mt���?      �?              �?      �?��RO�o�?              �?                       @       @                       @      �?      �?      �?ui��|��?�w�!�?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?      �?              �?m+�oM�?�?Y�?                      �?      �?      �?      �?       @      �?       @       @       @       @               @       @              �?�����f�?��x^�5�?      �?              �?        ��.�d��?      �?       @      �?       @               @       @                       @      �?      �?!����Z�?�e�\��?                                �'�K=�?      �?       @      �?                       @               @       @              �?      �?�Τ=���?��%���?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?E�(Ţe�?Z�ߜ�u�?                      �?        F���@��?              �?                               @               @       @              �?        �I�:Bl�?(��@�'�?                      �?      �?!�
���?      �?                       @       @       @       @       @       @       @              �?%K!�i�?��Z#PB�?              �?                �V�H�?      �?       @      �?               @       @               @       @              �?       @z�D_r�?���
��?                      �?        H���@��?      �?              �?               @       @               @       @                       @	{�����?�ީ�`|�?                                ��RO�o�?      �?                               @                                                       @�%��f��?�X�|�?                      �?        ���.�d�?      �?                               @       @       @               @       @      �?      @�Y e��?�I���?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      �?E�(Ţe�?�<��^?      �?                        ���V،?      �?       @      �?       @                                       @                      @,u�ئ�?��eHqm�?                      �?      �?�
��V�?      �?       @               @       @               @       @              �?      �?      �?�N���?��X	I��?      �?              �?      �?6���?      �?       @               @       @       @       @                       @              �?AIE���?Sm\2�?      �?      �?      �?        ?���@��?              �?                               @                                      �?       @�\d����?��.骀�?      �?                        	��V��?      �?       @      �?                       @       @                      �?               @3���?�`>�^��?      �?                      �?��RO�o�?      �?                       @       @       @       @               @       @                �cX�~k�?j�S߬��?      �?                        e�v�'��?      �?                       @       @                       @               @      �?        o��R��?�:�E���?      �?      �?                ���Vج?      �?       @      �?               @                               @              �?       @�hY7��?��8�g��?      �?              �?        �]�����?      �?                                                       @              �?      �?      @�Gm?C�?l^)s.��?      �?              �?        �@�6�?      �?                                                                              �?        ���G���?��`�P��?                                              �?              �?                                                              �?      @���S��?]�ׇx?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @$�$0�	�?����d1?      �?                                      �?       @                               @                                               @��ǰ2��?�\[L��p?      �?              �?        �@�6�?      �?       @      �?                                                              �?       @S,ZV��?���ַ?              �?                ���Vج?      �?       @      �?                                       @                      �?      �?S,?(��?7�09>�?      �?                                      �?                                                                                      @+�����?�'����i?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?tf�r��?      �?              �?      �?              �?              �?                                               @              �?       @O�)���?1~c�-l}?                      �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�d�Q�ϐ?t?Fg\�?      �?              �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?                �X����? zG�*�?                                �'�K=�?      �?       @               @                                       @              �?        ���Z��?n��	Ӽ?                                �'�K=�?      �?                       @                       @               @                        MaJ̖p�?ǜ��pj�?              �?                      �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?��9���?�:?y�?      �?              �?      �?P�o�z2�?      �?       @      �?       @       @       @       @       @       @       @      �?        C؋�ߵ�?J�����?      �?      �?      �?        3~�ԓ��?      �?       @      �?                                                              �?       @�ae��	�?`j��/��?      �?                        e�v�'��?      �?              �?       @               @       @                      �?               @a�:�?�`�1}�?      �?      �?                �K=��?      �?              �?       @       @               @       @       @       @      �?       @)���G��?��J�i�?                      �?      �?3~�ԓ��?      �?                       @                                               @      �?        �{B���?�����?      �?              �?      �?��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��w����?寚��?      �?              �?              �?      �?       @      �?               @       @               @       @       @      �?        7��+	�?<������?      �?                        �z2~���?      �?       @      �?               @       @       @       @       @              �?      @�U:'�?'����,�?      �?      �?      �?        �z2~���?      �?       @      �?               @       @       @       @              �?      �?        ]d�����?@�2�{��?      �?      �?                ��Vؼ?      �?       @      �?                       @               @       @              �?       @����e0�?�.�/���?                                              �?                                       @       @       @       @      �?              �?]�;x��?j�v<#z?                                �RO�o��?      �?       @               @               @       @                      �?               @�1����?)��=���?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?Y=4���?      �?      �?      �?        F���@��?      �?       @      �?                       @               @       @              �?       @�ߵN���?�+5�%�?      �?                        �]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�X����?|�5~�٧?                      �?      �?�K=��?      �?       @      �?                       @       @       @       @       @      �?        O|x�/��?��E����?      �?                        ��.�d��?      �?              �?                       @                       @              �?      �?:]��#��?UW�~n��?      �?                        �D+l$�?      �?              �?                                       @       @              �?       @���@���?1����5�?                      �?      �?P�o�z2�?              �?                       @       @       @       @       @       @              �?�5\.2��?|���4�?              �?                e�v�'��?      �?       @                       @               @       @              �?              @���q%�?X&s��?                      �?      �?��Vؼ?      �?              �?                               @                              �?       @
n��W�?kt����?      �?                        ���@��?      �?       @                               @       @               @       @                >�/�Q�?�����?      �?      �?      �?        Zas �
�?      �?       @      �?               @               @                      �?      �?        �}�m�?�B�ҹR�?      �?              �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ��Po��?��]�J�?      �?      �?      �?        6���?      �?       @      �?       @       @       @               @       @      �?      �?       @-����?a�n�%�?      �?                        $Zas �?      �?              �?                       @       @                      �?               @EDDDDD�?��v���?      �?              �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?                      @ś�8j��?���4�:�?      �?              �?      �?{2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?���sW�?                      �?      �?      �?      �?       @               @       @       @       @       @       @       @              �?9�WH�%�?VΊ��~�?      �?                        ?���@��?      �?                                                                                      @�9�፿�?���ܗ?      �?                                      �?              �?                                       @       @              �?       @ J�hY�?���f��?                      �?      �?      �?              �?                       @               @       @       @       @              �?B����?w��k���?                                �'�K=�?              �?               @       @               @                      �?              �?�w����?0�k�n�?      �?                        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @^��Z��?�qPh��?      �?              �?      �?F���@��?      �?              �?                       @               @       @                       @rv��?v���n�?      �?              �?        !�
���?      �?                       @       @       @       @       @       @       @      �?      �?ئ�N��?ط����?      �?      �?      �?        [as �
�?      �?       @      �?       @                               @                               @[ݧ����?R����?      �?              �?      �?P�o�z2�?      �?                       @       @               @       @       @       @                �Po���?݊�B�?      �?              �?        �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�d�Q�ϰ?� �'w�?                                �'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?���6�?fc≋�?                      �?      �?      �?      �?       @               @       @       @               @       @       @      �?      �?.2�z���?��CJ���?      �?                        �o�z2~�?      �?       @               @       @       @       @                       @                �A6w\I�?c8�S�'�?      �?                        6��9�?      �?       @               @                                                      �?      �?,u�ئ�?^��A�:�?      �?              �?              �?              �?               @       @       @                               @                B6w\I`�?hJ7o��?                                Zas �
�?      �?       @                       @       @       @       @       @       @              �?*1[�yj�?a|��l��?      �?                                      �?              �?                               @                                       @�/�Q��?d��"z?      �?              �?      �?              �?              �?                                                              �?       @������?B֜�#�x?      �?              �?      �?�z2~���?      �?       @               @       @               @       @               @              �?��Po��?v��S���?      �?              �?      �?              �?              �?               @                                                      �?����9��?��P�_z?              �?                �ԓ�ۥ�?      �?       @      �?       @                               @       @              �?       @��?y4��?t�1���?      �?                        �@�6�?      �?                               @                       @                               @H���<�?Ck�M�?                      �?      �?�'�K=�?      �?              �?               @                       @       @      �?      �?       @���`p�?4�yD=_�?                                ���Vج?      �?              �?                                       @                      �?      �?�����?T(j�K�?                      �?        �D+l$�?      �?              �?       @               @                              �?      �?      �?\�՘H�?'ڢ��?              �?                �
��V�?      �?       @      �?                       @               @       @      �?      �?       @w\I`��?�Xu��?                                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                        ]����`�?� �°�?                                �
��V�?      �?              �?                                               @              �?       @r�g�L��?��S�p�?                      �?      �?��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �k�.M��?�:'���?      �?                        �z2~���?      �?       @      �?                       @       @       @                      �?      �?��!�
�?��+r��?      �?                        ���V؜?      �?              �?                       @                       @                      �?1v�z�?v�:��?      �?              �?      �?���V،?      �?                                                                              �?       @K�*g��?���y�ր?      �?      �?      �?        ,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?,1[�yj�?{B��y�?                                �z2~���?      �?       @      �?               @                       @       @              �?      �?]d�����?P���x�?                      �?      �?��V��?      �?       @                       @               @       @       @       @      �?        )�tN|x�?�����?                      �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?��?��?                                F���@��?      �?                                               @       @                      �?      @��¯�D�?8��"�v�?                      �?      �?���.�d�?      �?       @               @       @       @       @       @       @       @      �?      @���l	�?Z��{i�?      �?              �?      �?	��V��?      �?              �?                                                              �?       @�돗�(�?O\���?                      �?        �z2~���?      �?                               @                                              �?       @~5&��?q���Ɇ�?                                �@�6�?      �?       @      �?                                       @       @              �?        ������?=%O���?                      �?                      �?                                                                              �?       @�{'Y��?���V�h?      �?                        6��9�?      �?                       @                       @       @                                s��2�?��#n7��?      �?              �?        !�
���?      �?       @                                       @       @       @       @      �?        """"""�?�.�/��?                      �?      �?�ԓ�ۥ�?      �?       @      �?               @       @               @       @              �?       @e����I�?ʑ�m�?      �?                      �?�D+l$�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ��C��?"!+��ϴ?      �?              �?        SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?       @               @�����`�?˟< �?                                [as �
�?      �?       @      �?                       @                       @              �?       @8�B�]��?w1�3��?                                SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����'t�?��.uc��?      �?                                      �?                                                                              �?        �bѲ
n�?�R�q�g?      �?              �?        >�]���?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?8�]�FR�?>:_e]�?                      �?      �?�K=��?      �?                       @       @       @       @       @       @       @              @�iŽ�,�?������?                                ���V؜?      �?                                       @               @       @      �?      �?       @��j1v�?G�0��ӗ?                                ���V،?      �?       @      �?                                       @       @              �?       @?(�tN|�?ў:?y�?      �?              �?        �ԓ�ۥ�?      �?       @      �?                                       @       @              �?       @c9�W�?���i��?      �?                        3~�ԓ��?      �?                                                       @       @      �?      �?        �\d����?��;Ͼl�?                      �?      �?3~�ԓ��?      �?                       @       @       @       @                       @              @-����?F��(���?                      �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?n��W�?A����z�?                      �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @����[�?�R�qޗ?      �?              �?        �@�6�?      �?       @      �?                                                              �?       @���I�:�?��VĨ?      �?                      �?p�z2~��?              �?               @                       @                       @              @۴��I�?�^���?                      �?      �?���.�d�?      �?       @      �?       @                       @       @       @      �?      �?        A���Kn�?��|!.��?                      �?      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?�ͪ�!��?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?"ApdL_�?      �?              �?      �?��.�d��?      �?                               @       @       @       @              �?      �?       @����`�?w�5(��?      �?      �?                v�'�K�?      �?       @      �?               @       @       @       @       @      �?              �?V�ߚ ��?i�$d�_�?                      �?      �?ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?       @                ����'t�?.!P��?      �?                        6��9�?      �?              �?                               @               @      �?      �?      �?�$0�	�?�L�p7�?                                $Zas �?      �?                                               @               @      �?               @���+$�?�7J-�?              �?                �z2~���?      �?              �?       @                                                      �?        /M��o2�?ПK ���?              �?      �?        $Zas �?      �?       @      �?                               @       @       @              �?       @;�RG�m�?�.B��?      �?              �?        p�z2~��?      �?       @      �?                       @               @       @              �?       @/��:]�?�X�i��?                                ���Vج?      �?       @      �?                       @       @                              �?       @9��_���?r����?                                �'�K=�?      �?                       @                               @                      �?       @ٴ��I��?�8fʹ�?                                �
��V�?      �?       @      �?               @                               @              �?       @��7q��?"���V@�?      �?              �?                      �?              �?                                                              �?       @�Kn��4�?��J�w?      �?              �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @���C�?��5b��?      �?                        �z2~���?      �?       @      �?                                       @       @              �?       @�i����?kj����?                      �?        ,l$Za�?      �?                       @       @       @                              �?      �?      @�:Blӊ�?�.��?                                ��.�d��?      �?       @               @               @       @       @              �?              �?�/�Q��?;h����?                      �?      �?              �?              �?               @                                              �?       @�6��`��?5� ��kz?      �?              �?              �?      �?       @      �?       @       @       @       @               @       @                ������?��>���?      �?              �?        !�
���?              �?                       @                                              �?      �?_W-��?{�$AP�?              �?      �?        v�'�K�?      �?       @      �?                       @       @       @       @      �?      �?      �?�<5���?"_m����?      �?                                      �?       @      �?                                       @                               @�s��2�?+T�ʟ?              �?      �?         �
���?      �?              �?                       @               @                      �?      �?1v�z�?�j,��@�?      �?                        �D+l$�?      �?                       @               @                               @      �?      @;�^!��?l�ZNy&�?      �?              �?      �?���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @E�(Ţe�?��Ki�.�?      �?                        6��9�?      �?              �?       @               @               @       @      �?      �?       @i�ae���?���o�?                                (�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?      �?WH�%���?��Yķ�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                        n��W�?�^/��"?                      �?      �?F���@��?      �?       @                                                                               @d��ht�?���S��?      �?                        6���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �m��W�?��m��?      �?                        >�]���?      �?       @      �?               @               @               @              �?       @�Gm?C�?��ч��?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @^��Z��?L�o#�V�?                                ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�X����?�[,�{�?      �?                                      �?       @      �?                                                              �?       @���6�?��H���z?                      �?        6��9�?      �?       @      �?                                       @                      �?       @�������?��%�>��?                      �?      �?�K=��?      �?       @      �?       @                       @               @      �?      �?      �?|]�;�?I��X�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                       @�d�Q�ϐ?���2�>r?      �?              �?      �?	��V��?      �?       @               @                       @                      �?      �?      @�<5���?���)׿?                                �z2~���?      �?       @      �?                       @               @       @              �?        w\I`��?��la��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @1[�yj�?؄�3��(?      �?                        ܥ���.�?      �?       @      �?               @       @               @       @       @      �?        �KS}��?������?                                3~�ԓ��?      �?              �?                       @       @       @              �?      �?      �?�^!ї��?p�i�?                                �
��V�?      �?                       @                                                      �?      �?�Po���?�
����?      �?                        �'�K=�?      �?                                                                                      @T�����?��^����?              �?      �?        �@�6�?      �?       @      �?                       @       @       @       @              �?        �#�d�Q�?w��|w�?                      �?      �??���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @9�%��}�?ӽ���t?      �?                        p�z2~��?      �?                               @                                              �?      @�b��!�?;E��`��?                                �D+l$�?      �?              �?                               @       @       @      �?      �?        �FR,?�?��(X�?      �?                        F���@��?      �?              �?                                                                        �Kn��4�?"��i«?                      �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @Y�)L�ْ?���Z�E�?              �?      �?        �@�6�?      �?       @                       @       @                       @      �?                Ȱ2���?mG�Z���?                      �?      �?!�
���?      �?       @      �?       @       @                               @              �?       @����C�?��ʪJ��?      �?                        ��RO�o�?              �?               @       @                               @              �?        +�����?6^�����?                      �?      �?�]�����?      �?                               @                                                      @:�X�?P5`����?                                              �?               @      �?      �?      �?      �?      �?      �?                        �d�Q�ϐ?�9�(� ?                                �ԓ�ۥ�?      �?       @                                                                      �?       @ e��h�?iR!|�l�?                      �?      �?�K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�?G���ܹ?                      �?      �?��.�d��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�X����?�UAZ�?                      �?      �?�K=��?              �?               @       @                                       @                t3NaJ��?�q2s��?                      �?      �?F���@��?      �?                       @                                                              @Q,?(��?m@r[���?      �?                      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              @F��1��?����S�?      �?              �?      �?,l$Za�?              �?               @       @       @       @               @       @      �?      �?t3NaJ��?�e5�g�?              �?      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?        ���̱�?@[W��?      �?      �?                F���@��?      �?       @      �?                                       @                      �?       @y4��0�?+�-L14�?                      �?        ��ۥ���?      �?       @      �?               @       @               @       @       @      �?        ���Kn��?6����?      �?              �?        v�'�K�?              �?               @       @       @       @       @               @      �?        2��l�?zb2X��?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                      �?F��1��?k�7�O�?                                �z2~���?      �?       @      �?                               @                              �?      �?q
Sb���?b��څ��?                                �]�����?      �?       @      �?                               @       @                      �?       @��,u���?%e���+�?                                F���@��?      �?              �?                                       @                      �?       @�j1v��?�����?              �?      �?        �K=��?      �?       @      �?       @       @                       @       @      �?      �?       @������?|>XT^1�?      �?                        ���V؜?      �?                               @                                              �?      @���'�?�����M�?                                ?���@��?      �?       @      �?                                                              �?       @�B�]�F�?�$1!���?                      �?      �?      �?      �?       @               @               @       @       @       @       @      �?      �?>�� Q��?�/׽~�?      �?              �?      �?�ԓ�ۥ�?      �?              �?               @               @       @               @      �?      @��J�ć�?c�KI���?      �?      �?      �?        6��9�?      �?              �?                                                              �?        *g��1�?�Y�̞��?      �?              �?                              �?                               @               @       @              �?       @���7q�?�?���m?                                F���@��?      �?              �?                                                              �?      @X-�r�?�T>E�?                      �?        ���@��?      �?       @                               @               @       @      �?                ����J�?[:���|�?      �?              �?      �?e�v�'��?      �?       @               @       @               @                       @      �?      �?��a/�?�L9�3�?              �?                ���V،?      �?              �?                                               @              �?       @4�G�Ɉ�?�"���Ӕ?      �?                      �?>�]���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�^W-��?������?      �?      �?                �@�6�?      �?       @      �?                       @               @       @              �?       @ʣ��8��?�s�����?                                �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @O�)���?&K(�%��?      �?                        �z2~���?      �?                       @               @               @       @              �?       @�z�D_�?�����	�?      �?                      �?p�z2~��?      �?                       @       @                                              �?       @��W��?-z�8v�?      �?              �?      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?                �����`�?�;�]��?      �?                        �
��V�?      �?       @      �?       @       @                               @              �?      �?V�;�RG�?��06V��?      �?                        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @Rp�l?�H�v�?      �?                      �?6��9�?              �?                                                                      �?      �?��C��?����*�?                              �??���@��?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @n��W�?Fy�S�~?      �?              �?        H���@��?              �?                       @                       @       @       @              �?O�)���?E�]���?              �?      �?        ��RO�o�?      �?              �?               @       @       @       @              �?      �?       @��1��?�|�:��?      �?              �?      �?��ۥ���?      �?                       @               @       @               @       @      �?      �?�9�፿�?��ÙK�?      �?              �?      �?      �?      �?                       @       @               @       @               @                ��,����?�c���?      �?                        ���V؜?      �?                                       @                                      �?       @���w��?O�\���?      �?              �?        v�'�K�?      �?       @               @       @       @                               @      �?      �?��3��x�?��uH�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @M:'>��?b:���9+?      �?      �?      �?        �@�6�?      �?       @      �?                       @                                      �?       @�:]���?#�Uj9�?                                ���V،?      �?              �?                                       @                      �?       @~5&���?b�/
b7�?              �?                ��RO�o�?      �?       @      �?               @                                              �?       @L���S�?6̾�|��?      �?      �?                ���Vج?      �?              �?                                       @       @              �?       @���¯�? d����?                      �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?m+�oM�?W@z�y�?      �?              �?        Zas �
�?      �?       @      �?               @       @       @       @       @              �?       @W����?�E�HFD�?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        ��?y4��?zNN�c��?              �?      �?        �
��V�?      �?       @      �?               @       @       @                                       @��ǰ2��?濐f��?                      �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @#w\I`ޓ?Z䣒�{�?      �?              �?      �?�V�H�?      �?       @      �?               @                                              �?        M+�d��?�+mIz��?                      �?        p�z2~��?      �?       @      �?                                                              �?      �?/M��o2�?E 5p��?                                              �?       @      �?                                               @              �?       @�_���@�?lߤJ?              �?      �?        ��V��?      �?              �?               @       @       @       @       @       @      �?      �?[�KS}��?������?                      �?      �?��ۥ���?      �?       @      �?       @       @       @       @       @       @       @                �B�/���?���?l��?      �?              �?        [as �
�?      �?       @      �?                       @               @                              �?*1[�yj�?MIDMU��?              �?                Zas �
�?      �?                                               @       @                               @���?y4�?�2�
���?                      �?        6���?      �?       @      �?       @       @       @               @       @       @      �?        :�$0�	�?�%�\���?                      �?      �?��.�d��?      �?              �?       @               @       @                              �?        
Sb����?�m����?      �?                        �o�z2~�?              �?               @       @       @       @                       @      �?        �Kn��4�?ƿZ �2�?                                ��Vؼ?      �?       @      �?                                                              �?      �?""""""�?�e�qE+�?                      �?      �?3~�ԓ��?      �?       @      �?               @                       @       @              �?       @��l	��?
����?                      �?        ���V،?              �?                                                       @              �?       @l��4�u�?�k�q�w?      �?                                      �?              �?                                                              �?       @X-�r�?�3�
'x?                                �'�K=�?      �?       @      �?                                       @                      �?       @���C��?�`�'��?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @nC��x�?�|�:�?              �?                �@�6�?      �?       @      �?                                       @       @              �?        r@���?�y��?��?                      �?        ��Vؼ?      �?              �?                                       @       @                       @[ݧ����?cmweU��?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @\��r�?�:u߁�?                                ���Vج?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?�U�����?��B.�O�?      �?                         �
���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�፿Po�?�I��?      �?      �?                ��V��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        �j1v�?鐷�@}�?              �?      �?        �z2~���?      �?       @      �?               @       @               @                      �?       @7���l�?�j4,�þ?      �?      �?                F���@��?      �?                               @                       @                      �?       @Ήo���?.�����?                      �?      �?���V،?      �?              �?               @                                              �?        ���G���?�|�:�?      �?                        ���V،?      �?              �?                       @               @       @                       @3��l�?o�vo�Ғ?              �?                F���@��?      �?              �?       @                                                                0�	��?��Ĳ���?      �?                        ���Vج?      �?              �?                               @       @       @              �?       @�4�G���?�:�&C��?      �?              �?      �?$Zas �?      �?       @      �?                       @               @       @      �?               @.�jL��?�"b�/�?                      �?        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                b��1��?9]n���?      �?              �?        �ԓ�ۥ�?              �?               @               @               @       @      �?              �?��r�9�?
U&>�?                                 �
���?              �?                               @       @       @                      �?      �?�r@��?���>5�?      �?              �?      �?3~�ԓ��?              �?                               @               @       @                      �?F�X�ڙ�?�a�$�?                                              �?              �?       @       @               @                              �?      @"�
���?�E���~?      �?                        �@�6�?              �?                       @               @                              �?      @L��b��?����}�?                                �
��V�?              �?                               @       @                              �?      @۴��I�?zb2Xػ?                      �?      �?6��9�?      �?                               @       @                                      �?      @.������?JBV�u�?              �?      �?        >�]���?      �?       @               @       @       @       @                      �?      �?      �?yjH���?TS�[Z��?                              �??���@��?              �?               @       @       @               @       @              �?      @~�ɣ���?wB ��7�?      �?              �?        p�z2~��?      �?       @      �?               @       @               @       @              �?       @�X����?\���:��?                      �?        p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����[�?���lq�?              �?                              �?              �?                                       @       @              �?       @�+	�{B�?\��J5"�?                      �?        ���V،?      �?       @      �?                                       @                      �?       @
Sb����?��&��<�?                      �?      �?��V��?      �?              �?                       @               @       @      �?      �?       @����C�?j�w���?                                ���V،?      �?              �?                                                              �?       @���S��?+u-Ye�?              �?                              �?              �?                       @                       @              �?       @�_���@�?lߤJ?      �?                        ,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?nC��x�?˟< �?      �?                        >�]���?      �?       @      �?               @                       @       @                       @�Τ=���?굽���?                                �ԓ�ۥ�?      �?       @      �?                       @               @       @              �?       @��2�?�R���?                                �'�K=�?      �?                       @                       @                      �?                ���@���?�L���W�?      �?                        e�v�'��?              �?               @       @                               @       @                 �����?��&vQ��?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?                      @����'tx?�C���?      �?                      �?��.�d��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�U�����?�\��޺?      �?              �?      �?��RO�o�?      �?                       @       @                       @                      �?       @_W-��?�f�[$�?      �?      �?      �?        6��9�?      �?       @      �?                                               @                       @�}�m�?�O?���?      �?              �?        6���?      �?                       @       @       @                              �?              �?�5\.2��?��3.�?                      �?      �?�K=��?      �?       @               @                               @       @       @      �?       @���I�:�?�EF�=�?                                �@�6�?              �?                                       @       @       @      �?      �?      @!�iŽ�?L!>�!��?      �?              �?      �?$Zas �?      �?              �?               @                       @                      �?      @V�i���?�*��-��?                      �?      �?�]�����?              �?               @               @       @       @       @      �?      �?      �?a/���?60�\�?                                Zas �
�?      �?       @      �?                       @                       @                      @��ߵN��?�A���=�?              �?                �z2~���?      �?       @               @                       @               @              �?       @���"X~�?dA"�Xz�?      �?                        �V�H�?      �?                                                                              �?      �?���8�)�?V۾�9�?              �?      �?         �
���?      �?       @      �?                       @               @       @              �?        7���l�?�	4g�?      �?              �?        >�]���?              �?                               @       @       @       @      �?      �?        t3NaJ��?���lF��?      �?                        �@�6�?      �?       @                               @                       @      �?              @I!�i��?忐f��?              �?                ���V؜?      �?              �?                                                              �?       @�V�ߚ�?4.��k��?              �?      �?        �]�����?      �?       @      �?       @               @       @       @       @      �?      �?      @�C��?���G��?      �?                      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?                        #w\I`ޓ?�V�φn?      �?                        ���Vج?      �?                                       @       @       @       @                        _W-��?��.em�?      �?              �?        ��ۥ���?      �?       @      �?       @               @       @       @       @       @      �?      �?�l��?���ݨ�?      �?              �?      �?      �?      �?       @               @               @       @                       @      �?      �?��C��?c�񉦲�?      �?              �?        �RO�o��?      �?       @      �?                       @               @       @       @              �?�3i�ae�?�,�=�U�?                                �z2~���?      �?                                                                              �?        �{'Y��?rD��^ޭ?      �?      �?                              �?       @      �?                                                              �?       @0�	��?�^�?{?      �?              �?      �?P�o�z2�?      �?       @               @       @       @       @       @       @       @      �?      �?Gm?C؋�?G��ci��?      �?                        ���Vج?      �?       @      �?               @       @                       @                       @�Up�l��?%��ӗo�?                      �?      �?$Zas �?      �?       @      �?                       @       @               @              �?        ��[�՘�?�%'�y�?                      �?        ���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?)g��1�?		#�a!�?      �?              �?      �?��Vؼ?      �?                               @               @                                      @R��'�F�?b�/��?      �?      �?      �?        3~�ԓ��?      �?       @      �?                                               @                       @ J�hY�?�� ���?              �?      �?        ,l$Za�?      �?       @      �?                       @       @       @       @                       @q���Y�?Q6^���?                      �?      �?�
��V�?      �?       @      �?       @       @                                              �?       @�vAI�?�8�����?                              �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?nC��x�?_�;[w��?      �?              �?      �?��ۥ���?      �?       @      �?       @               @               @       @       @               @��+	��?�:Z�F�?      �?      �?      �?      �?�K=��?      �?       @      �?               @       @       @       @       @              �?       @���<��?� ,�H��?              �?                ���V،?              �?                                                                               @��*��?�R��e?      �?                        �'�K=�?      �?                                       @       @       @       @      �?      �?        k� 6\.�?�(!�n�?      �?                        p�z2~��?      �?                       @                       @                                       @䶺O_�?��,S��?                                �ԓ�ۥ�?      �?       @      �?                                       @                      �?       @��`�AQ�?3(�����?              �?      �?      �?�K=��?      �?       @      �?               @                                              �?      @4�G�Ɉ�?�	1����?      �?                        F���@��?      �?       @      �?                                       @       @                       @Aʾ����?����W�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?n��W�?�o�ݙ?      �?              �?        v�'�K�?      �?       @      �?       @       @       @       @       @       @      �?                E�Ή�?���i�A�?                                �@�6�?      �?                       @               @       @       @       @      �?      �?        ��*��?Ys��b�?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        ��ht3�?K%,h�c�?                      �?        Zas �
�?      �?       @      �?                               @       @       @      �?                �3i�ae�?�����?                                ��ۥ���?      �?       @      �?               @                       @       @              �?       @9�)1[��?��"��?                      �?      �?e�v�'��?      �?       @                       @       @       @       @       @              �?       @�a�(Ţ�?�o;Ԣ�?      �?                      �?6��9�?      �?       @      �?                                       @       @                       @��a��?�����?      �?      �?      �?        �
��V�?      �?       @      �?                                                              �?       @�/�Q��?I	.����?                                �@�6�?      �?              �?                       @       @               @              �?       @O��b��?{Ν�6��?      �?              �?        H���@��?      �?       @                               @                                              �?.������?�W3�z�?      �?                                      �?              �?                                       @       @              �?       @�p��R�?�ѐ �o�?      �?      �?                �6��?      �?                               @       @       @       @              �?      �?      �?'#��~��?��x��M�?      �?              �?      �?���V،?      �?                       @       @               @                       @              @��¯�D�?H���e�?      �?                                      �?              �?                                               @              �?       @�:]���?8rK��M}?                                �D+l$�?      �?                       @                                                      �?      @d��ht�?��J��k�?      �?      �?      �?        �]�����?      �?              �?               @       @               @       @      �?      �?        ���?y4�?)H���?      �?              �?        ��Vؼ?      �?              �?               @       @       @       @                      �?      @�g�L�c�?(�8����?      �?              �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?m+�oM�?��z�o�?                      �?        �@�6�?      �?       @      �?                                       @       @              �?       @J�hY7�?i�_�
��?                                ?���@��?      �?                                                                              �?      @*g���?�DkJ���?      �?                        ���V؜?      �?              �?       @                       @                              �?      @]��#�d�?�m_���?      �?              �?        (�K=�?      �?       @                       @       @       @       @               @              �?�cX�~k�?U�Oˊ^�?                      �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�d�Q�ϐ?ms��?      �?                        ?���@��?      �?       @      �?                                                              �?       @�c=kg�?8 X���?                      �?      �?p�z2~��?      �?       @               @       @               @       @       @       @      �?      �? J�hY�?1x��1�?                              �?	��V��?      �?       @      �?               @       @       @                              �?      �?�X�ڙ��?'�3���?      �?      �?      �?        �'�K=�?      �?       @      �?               @                               @              �?       @t3NaJ��?d���-�?                      �?      �?���Vج?              �?                       @               @                                       @�����`�?^�XO��?      �?              �?        �RO�o��?      �?              �?               @                       @       @      �?      �?       @�FR,?�?������?                      �?        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?m+�oM�?��u��?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              @����'t�?���`Q�?                                	��V��?      �?       @      �?                       @                                                ���w��?�4���?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ,1[�yj�?�t�c���?                      �?        ���V،?      �?              �?               @       @                                                �j1v��?B�� �F�?      �?              �?      �?��RO�o�?      �?              �?       @       @                                      �?      �?      �?7w\I`��?ھ�9.�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @-h#���?�T����?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @m+�oM�?`�I���?                                 �
���?      �?              �?                                       @       @              �?        r�9ֳv�?����[��?      �?      �?      �?      �?�RO�o��?      �?       @      �?       @       @                               @              �?       @HT�n��?]k7�@�?                                F���@��?      �?       @      �?               @                                              �?        333333�?]o/2ɭ?                      �?      �?�V�H�?              �?               @       @                                                        ^�(Ţe�?����l��?                                ���V،?      �?              �?                                                              �?       @'#��~��?a��}pЈ?              �?                >�]���?      �?       @               @               @       @               @       @                h>�/��?ѽ@�Z��?      �?      �?      �?        	��V��?      �?       @      �?                                       @       @              �?       @����_�?�6T�Z��?      �?                        �@�6�?              �?               @                       @       @                      �?      @T�����?��/�8S�?      �?              �?      �?p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ò
n�ͭ?I)�˰?                      �?      �?�o�z2~�?      �?                       @               @       @       @              �?      �?        L�*g��?Y8��X�?      �?              �?        (�K=�?      �?              �?       @       @               @                       @                l	�Y �?����Q �?      �?              �?      �?$Zas �?      �?              �?                                                              �?       @��J��?�d��r�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @��N�ԑ?߃�U�Җ?      �?              �?      �?��RO�o�?      �?       @               @       @                               @                      @�c9�?�ȍ��Y�?              �?      �?        	��V��?      �?       @      �?       @               @                                      �?        ��>|]�?�H݇V�?      �?              �?      �?>�]���?      �?       @      �?                       @       @       @       @       @      �?       @���I{�?e�5c���?      �?              �?      �?F���@��?      �?                       @                                                      �?      @uN|x�/�?8v��_̰?      �?                        6��9�?      �?                               @                       @                      �?      @.��:]�?[@��Q�?      �?                        ��Vؼ?      �?       @      �?               @                       @       @              �?      �?��E���?���Ε�?                      �?        SO�o�z�?      �?       @       @      �?      �?      �?      �?      �?      �?       @               @��N�Ա?H|�$A�?                                ���V،?      �?       @                       @                                                      @^!ї��?�r�`��?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @              @E�(Ţe�?��`���?                                �z2~���?      �?       @      �?               @                       @                      �?      �?}�mu��?ԛ�����?      �?              �?        ��ۥ���?      �?       @      �?       @       @       @       @       @       @       @      �?       @�e0
84�?�S-���?      �?                        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�0[�yjv?�1��ſ?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?               @       @       @       @       @       @      �?        ;�X��?,5�%��?      �?                      �?�@�6�?      �?                                                                                      @Z��r�?]� )2��?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?Y�)L�ْ?�XrS* ?      �?                        �z2~���?              �?               @               @       @                      �?                q����?�\��.��?                      �?      �?���V،?      �?                                                       @       @                      @�J�ć7�?5U�N�?      �?      �?      �?        F���@��?      �?       @      �?                       @               @       @              �?       @����?�\�u>�?      �?                              �?      �?       @      �?               @       @               @       @       @      �?        �=�� Q�?b�0TKy�?      �?                                              �?                                                                      �?       @b��1��?.�a���D?                              �?�K=��?      �?       @      �?               @               @       @       @      �?      �?        Ɉ���!�?١���?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                       @��1�~?���3�?                                6���?      �?              �?       @       @       @               @       @      �?      �?       @�(Ţe�? ����?      �?              �?        ��V��?      �?              �?                       @               @       @      �?      �?       @'t J��?�����I�?      �?                        �]�����?              �?                       @       @                       @      �?      �?        o�Wc"=�?��v<#�?      �?              �?        	��V��?      �?       @      �?               @                                              �?        �~5&��?��ɡx�?      �?              �?        ��Vؼ?      �?                                       @               @       @              �?      @���"X~�?R�φ�?                                �@�6�?      �?       @      �?                       @               @       @              �?        g�L�cX�?��Ī�?      �?                      �?H���@��?              �?               @                               @              �?      �?      �?�U�����?�{�m��?                      �?      �?SO�o�z�?      �?              �?                       @       @       @       @       @      �?       @GR,?(�?֢K����?      �?                        6��9�?      �?              �?                       @               @       @              �?       @p2��g�?�/@ȭm�?                                              �?               @      �?      �?      �?      �?      �?      �?                       @E�(Ţe�? ��??      �?              �?        �ԓ�ۥ�?      �?              �?                       @       @                                       @ݧ����?87�6�j�?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @      �?      @��%���?�{�� z�?                      �?        Zas �
�?      �?       @      �?                       @       @       @       @              �?       @����>�?��M��?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����'t�?54�Ǵ�?      �?              �?      �?p�z2~��?      �?       @                       @                                                       @���@���?9^��1��?      �?                                      �?                                       @                                      �?       @9��_���?fҫS�m?              �?                �@�6�?              �?               @                               @                      �?       @�*��?�F�C�?      �?      �?                ���V؜?      �?       @      �?                                                              �?       @�c=kg�?��E0+�?      �?      �?      �?        F���@��?      �?       @      �?       @       @                               @                      �?����C�?_��!Y�?      �?              �?        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�d�Q�ϐ?��?�?      �?                        ?���@��?      �?       @      �?                                                              �?        g��-�?"�Wi�?              �?                �ԓ�ۥ�?              �?                               @               @                      �?       @�X����?��Tq��?                      �?        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?                ���@��?R�3.z|?      �?              �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                )g��1�?t9��h�?                      �?      �?      �?      �?       @      �?       @       @       @               @       @       @              �?�C��?寚��?      �?      �?      �?        �K=��?      �?       @      �?               @               @       @       @       @                c��!��?�:J����?              �?              �?              �?              �?                                                              �?       @������?B֜�#�x?      �?                        �@�6�?      �?       @       @      �?      �?      �?      �?      �?      �?                      �?�Y;���?�D���?      �?                        �'�K=�?      �?              �?                       @               @       @              �?       @c9�W�?WSѭJP�?      �?                      �?�z2~���?      �?                               @               @                              �?        ��W��?<������?      �?      �?      �?        �RO�o��?      �?       @      �?               @       @               @       @      �?      �?       @}䛌8j�?w��V�?      �?              �?        (�K=�?      �?       @                       @       @       @       @               @                �}��j�?i�$d�_�?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�U�����?/Z0�-t�?                                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                      @�U�����?�g��?                              �?���@��?      �?                       @               @       @       @              �?      �?      �?o��z��?1�nE��?      �?                      �?�'�K=�?              �?               @                       @               @       @      �?      @�9�፿�?�J��H.�?                                ��RO�o�?      �?       @      �?                       @                                      �?       @*L����?oZ;���?      �?                        SO�o�z�?      �?       @      �?       @       @       @                       @      �?      �?       @�$K!��?3ң�"��?                                �z2~���?      �?                               @       @                              �?                ͤ=����?��P�U�?      �?                      �?                      �?                       @               @                                      @��<݌�?� >�!�[?                      �?      �?�]�����?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        h#���?�WQ�sȼ?              �?      �?        v�'�K�?              �?                       @       @               @              �?                O�0@�b�?�Z���7�?              �?      �?        ��V��?      �?              �?       @       @       @                       @                       @�FR,?�?eR�L��?      �?                        >�]���?      �?                               @               @       @       @      �?      �?        �ئ�N�?�����?      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @                �'�F7�?��	�j�?      �?              �?      �?�z2~���?      �?       @      �?               @       @       @       @       @       @      �?        �n�Wc"�?�m�n��?      �?              �?      �?�K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�%��f��?���a��?      �?              �?      �?>�]���?              �?                       @       @                              �?      �?      �?f{����?�]ݒ���?                      �?        P�o�z2�?      �?       @      �?       @       @       @       @       @       @       @              @��!����?u�w@o�?              �?                              �?       @      �?                                               @              �?       @H*��E�?	;�m,P?                                      �?      �?       @      �?               @       @       @       @       @       @      �?      �?�^!ї�?Rt����?              �?      �?        ��RO�o�?      �?       @      �?       @                       @       @       @              �?        ��0%f�?ͤe�>
�?                                                      �?                                                              �?              @����[�?��0�U�J?      �?                                      �?              �?                                                              �?       @ї�V�i�?:j)��x?      �?      �?      �?        �]�����?      �?       @      �?               @       @               @       @              �?       @���-��?��;�?                                ���V،?      �?                                       @                       @                       @Ƣe� �?Ye?�?                      �?        �V�H�?      �?       @      �?               @               @       @       @      �?      �?       @3��g�?�|�#���?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @              @^��Z��?�A@�QN�?      �?              �?      �?�D+l$�?      �?       @      �?               @               @                              �?        kg����?�u�ұ��?      �?      �?                              �?       @      �?                                                              �?       @k� 6\.�?_=?|�z?                                �@�6�?      �?       @               @               @       @               @              �?        �k�.M��?��8���?                                ���V،?      �?              �?                                                              �?       @Y�ڙ���?�2♁(�?              �?      �?      �?�V�H�?      �?       @      �?       @       @               @       @       @              �?       @��|�G�?�+_J�?      �?      �?      �?        �@�6�?      �?                       @       @                               @              �?        Ň7�B��?*�"����?      �?      �?                ���Vج?      �?                                       @                                               @���7q�?�ĪЙ?                                6��9�?              �?               @                                                              @eZq�$K�?���ع�?      �?                      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              @M:'>��?̈g��?                                �'�K=�?      �?                                       @       @               @                      @ٙ�ǰ2�?�2�V��?                      �?        �z2~���?      �?       @               @               @               @       @      �?               @���Z�K�?��\/X�?      �?              �?      �?      �?      �?       @      �?               @       @               @       @      �?      �?      �?z�D_r�?��:?y�?      �?              �?        ���@��?      �?       @      �?               @                       @       @      �?      �?       @�C��x�?��P�,��?                      �?      �?�z2~���?      �?       @      �?                                       @                      �?       @x�����?��K��?      �?              �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?����'t�?K@���?      �?      �?                              �?                                                                              �?      @ui��|��?b�S�	�i?      �?      �?      �?        �K=��?      �?       @      �?       @       @                                                        �'�F7��?ƈ)%W��?      �?                                      �?                                                                                      �? �����?�ꖜ��i?                      �?        	��V��?              �?                       @       @                                      �?      �?��D)�?�Jk���?      �?              �?        (�K=�?      �?                       @       @       @       @                       @              �?Ň7�B��?�����?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @-h#���?�>�]ݒ�?      �?              �?      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?\��r�?�l��?                      �?      �?���Vج?      �?              �?                               @       @                      �?       @�@��~�?(<����?                      �?      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�p�Ȭ?▿j�J�?      �?                                      �?              �?                                       @       @              �?       @R��'��?��4��?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?�9�(� ?      �?                        >�]���?      �?       @      �?       @                       @       @       @              �?      @�������?�v��S�?                      �?        6��9�?      �?                                                                                      @~PT���?s��q�?�?      �?              �?        !�
���?      �?                       @       @       @       @       @       @       @      �?      �?�'�F7��?0�h}��?      �?              �?      �?�@�6�?      �?       @      �?               @       @               @       @                       @A���Kn�?���s���?      �?      �?                ��ۥ���?      �?       @      �?       @                               @                      �?       @�
n���?&�P�@e�?                      �?      �?��ۥ���?      �?       @      �?       @       @       @               @               @      �?      �?�$K!��?�K.r��?      �?                        >�]���?      �?                       @               @                              �?              @Ln��4��?����)�?      �?                        �V�H�?      �?       @      �?               @       @       @       @       @       @               @	�p���?iX�=	�?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?               @       @               @              �?              �?d�#�6��?̳��U��?      �?              �?                      �?       @      �?                                                              �?        ����9��?��P�_z?      �?      �?                ���V،?      �?       @      �?                                                              �?      @̖p���?F��<\B�?              �?                ���Vج?              �?                                               @       @                       @��g{�?@Ր�,�?      �?              �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?\��r�?O9N�O,�?                      �?      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?}���p?                                (�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?2w\I`޳?g�[$�?                                      �?      �?       @      �?       @       @       @       @       @       @       @              �?�c=kg��?�����?      �?                        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @^��Z��?L]f�v�?      �?              �?        !�
���?      �?       @      �?               @                               @      �?      �?      �?����?q��`��?      �?              �?        ��V��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?���C�?� �P@��?      �?              �?        ���@��?              �?               @                       @       @              �?      �?        �r@��?�����?              �?      �?              �?      �?       @      �?       @       @       @               @       @       @      �?       @4i�ae��?�����?      �?      �?      �?      �?      �?      �?              �?       @               @       @       @       @       @      �?      �?�����U�?�c���n�?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @-h#���?+�TYx�?              �?                ���V؜?      �?       @      �?                                                              �?      �?��C��?zC��?                                �'�K=�?      �?       @               @                                       @              �?       @��3��x�?Y�RR)��?      �?      �?                �'�K=�?      �?       @      �?                       @                                      �?       @\�՘H�?�q����?      �?      �?                3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?-h#���?��{�Cΰ?      �?              �?      �?�z2~���?      �?       @                       @               @                       @              @�3i�ae�?A@�QN��?      �?              �?      �?      �?      �?       @      �?       @               @               @       @      �?      �?        )����?��Tq��?      �?              �?      �?P�o�z2�?      �?              �?       @       @       @               @       @       @      �?        5&����?N0k�?      �?                        �ԓ�ۥ�?      �?       @               @               @                                      �?       @��U�?GGp�-��?      �?      �?      �?        ��V��?      �?              �?       @       @               @               @      �?      �?       @������?uϋ�4m�?      �?      �?      �?      �?�'�K=�?      �?       @      �?                       @               @       @              �?       @e����I�?��f���?      �?              �?      �?6��9�?              �?               @       @       @       @               @       @              �?��Y;��?m�۳��?                      �?        	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @,1[�yj�?	���?      �?      �?      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      @6��w���?��Ds��?      �?                        H���@��?      �?       @               @       @       @       @               @                        ��e0
8�?՘�q=��?      �?              �?      �?��.�d��?      �?                       @       @       @               @       @       @               @��.h�?9�o����?                                ���V؜?      �?              �?                                       @                      �?       @)�tN|x�?�v�寚?      �?                        6��9�?      �?                                                                              �?      �?��j1v��?�����?                                              �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?@Ր�,?                      �?        �D+l$�?      �?       @                       @               @       @       @      �?      �?       @���U���?݊�B�?      �?                        �@�6�?      �?                               @                       @              �?      �?       @�N��b�?1#E�?      �?                        ��RO�o�?              �?                               @               @       @              �?       @ئ�N��?,�;c��?                      �?      �?�'�K=�?      �?              �?               @                       @                      �?       @kg����?a!�ʧ��?                      �?        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?                        ]����`�?P��<A�?      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?-h#���?87�6�j�?      �?                        F���@��?      �?       @      �?                               @       @       @                       @��¯�D�?��z���?      �?                                      �?                                               @                              �?       @���!���?UB����l?      �?      �?      �?              �?      �?       @      �?               @       @               @       @       @      �?        q���Y�?qm���S�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                nC��x�?8}����?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?�%�ۄ?              �?                ���V،?              �?                               @                                      �?       @���J�? �|��I|?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @#w\I`ޓ?g�&
�?      �?      �?      �?        �o�z2~�?      �?       @      �?               @                               @              �?        �hY7��?�'�ܷ�?      �?      �?      �?      �?�@�6�?      �?       @      �?                                                              �?      �?""""""�?��c�X�?      �?      �?                �'�K=�?      �?              �?               @                                              �?       @�u�b���?.)�$.�?      �?              �?      �?(�K=�?      �?       @      �?               @                       @       @       @                C�}�?ddМ�B�?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @,1[�yj�?^ųR	j?      �?                        �'�K=�?      �?       @                       @               @                              �?      �?,ZV���?��e=4�?      �?      �?      �?        �6��?              �?                                                                      �?       @�d�Q�ϰ?��杭�?      �?                        �]�����?      �?       @      �?               @                       @       @              �?       @H���<�?����?              �?      �?      �?              �?              �?                                                              �?       @o�Wc"=�?\��Kd�w?      �?              �?      �?3~�ԓ��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @��N�Ա?������?      �?      �?                �z2~���?              �?                               @       @               @              �?       @b����,�?�=	��?                                ��ۥ���?      �?       @               @               @       @       @       @      �?      �?      �?h{����?�3�e��?      �?                        e�v�'��?      �?       @      �?                       @                       @                      �?��%���?��4b��?      �?      �?      �?      �?Zas �
�?      �?       @      �?               @                       @       @      �?               @�$K!��?Gu[D��?                      �?        �D+l$�?      �?       @      �?                                               @              �?       @�_���@�?����=�?              �?                F���@��?      �?              �?                       @               @                      �?       @����?��Bt�?                                ���V؜?      �?       @                                               @                      �?       @z�rv��?PͿ���?                                              �?       @      �?                                       @       @              �?       @�q%�yO�?�e=4��?                                (�K=�?      �?       @      �?               @       @       @                      �?      �?        ���@���?�����?                      �?        �'�K=�?      �?       @                       @       @       @       @              �?                ����9��?"�B6�?                                SO�o�z�?      �?       @                               @       @       @       @       @      �?      �?��I{+�?ԓ��:��?                                	��V��?      �?       @      �?       @       @                       @                      �?       @�FR,?�?�Ru���?                      �?      �?ܥ���.�?      �?                       @       @       @                       @       @      �?      �?cX�~k��?!�����?      �?              �?              �?      �?       @               @       @       @       @       @       @       @      �?        ����!��?.o�C���?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�U�����?qpTV�?                      �?        ���.�d�?      �?       @               @       @       @       @               @       @      �?      @���[�??�4���?      �?                        ��RO�o�?              �?                               @       @       @       @              �?       @jL�*g�?B��~�?�?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�d�Q�ϐ?�*I��?      �?                      �?H���@��?      �?              �?               @                       @       @              �?       @�	�p��?]����?      �?                        �z2~���?      �?              �?                                       @                      �?       @h#���?āy��b�?      �?                        �z2~���?      �?                       @                       @                                      @����'t�?��ʲ?      �?      �?      �?        ��.�d��?      �?              �?       @               @       @       @       @      �?      �?        z�D_r�?v�K�+�?      �?                        ���V،?      �?                                                                                      @�d�Q���?��	�z?                                $Zas �?      �?               @      �?      �?      �?      �?      �?      �?              �?        nC��x�?Z�7J�?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����[�?�I�.�?      �?                        ?���@��?      �?       @      �?       @                                                      �?       @���U���?�G{߿�?                                �@�6�?              �?                                               @       @                      �?�{'Y��?rB�vr��?      �?                        �'�K=�?      �?       @      �?                                               @              �?       @&�1�L��?,a�����?      �?                        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @-h#���? 2���?      �?                        �'�K=�?              �?               @                                                      �?       @��*��?5/�CZ��?                      �?         �
���?              �?               @               @                              �?              �?�������?�IkZ�?                                ܥ���.�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?^Zq�$K�?�w�@G2�?                                ��RO�o�?      �?       @      �?               @       @               @       @       @               @��+	��?��Yԭ��?                                ��Vؼ?      �?                               @               @       @                              @f��1��?�q��Ʊ?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @              �?��O�n�?XC�#���?                      �?      �?���.�d�?      �?               @      �?      �?      �?      �?      �?      �?       @              @#w\I`ޓ?`�[��?      �?              �?        ���.�d�?      �?       @      �?               @               @       @       @       @      �?       @5&����?�C�~i �?                              �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?♁(�?      �?              �?        6��9�?      �?              �?                                       @                      �?       @�`�AQ��?��Vĸ?      �?              �?      �?      �?      �?       @      �?       @       @       @               @       @       @      �?      �?;�X��?������?              �?                �@�6�?              �?                                               @       @              �?       @?y4���?F1�}ܜ?      �?              �?        p�z2~��?      �?       @      �?                                       @       @              �?       @y���?WNڵ�v�?      �?                        6��9�?      �?                       @                                                      �?      @H*��E�?' ���?                                ���V،?      �?                               @                       @                      �?       @^��C��?�i����?      �?                      �?F���@��?      �?                                                       @       @                      �?�w�ӥ��?��0��?      �?      �?      �?        ��ۥ���?      �?       @      �?                                               @              �?       @�W���?�� W-�?      �?                        $Zas �?      �?       @      �?                       @               @                      �?       @��O�n�?'�U��?                                ���V،?      �?              �?                                       @                      �?       @7w\I`��?_I���?      �?                        ���V،?      �?                               @                                              �?      @ e��h�?#md��y�?                                SO�o�z�?      �?                       @       @               @               @      �?      �?      @��f��}�?�oC��%�?      �?                        6��9�?      �?                                                                                      @*g���?�z���?      �?              �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�X����?���3�?                      �?        �o�z2~�?      �?                       @               @       @       @       @       @              @�����?Y}��jW�?      �?      �?                ��RO�o�?      �?       @      �?                                       @       @              �?       @IE����?�Jk���?      �?                        �'�K=�?      �?       @      �?               @                       @       @                       @#s�g�L�?u�=7���?      �?                        H���@��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �k�.M��?;�ਬl�?                                p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����`�?��}U�ݽ?      �?      �?      �?        �z2~���?      �?       @      �?               @       @               @       @              �?       @z�D_r�?��vgL��?                      �?      �??���@��?      �?              �?                                               @                       @B�/����?��5�Ơ?      �?      �?      �?        ��RO�o�?      �?       @                       @       @       @       @       @              �?        y4��0�?û.m���?      �?                        �'�K=�?      �?                       @               @               @       @       @      �?        ,�����?�9�[޾�?                                �'�K=�?      �?       @                       @                                      �?      �?       @
84���?�p�j<��?                                F���@��?      �?                       @                               @       @              �?       @����7�?`�`��?                                	��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�፿Po�?U�y�?                      �?      �?Zas �
�?      �?              �?               @                                                        h>�/��?��)�Lb�?                                �@�6�?      �?                                       @       @                      �?                �G�Ɉ��?.�KQ ��?              �?      �?      �?��V��?      �?       @      �?               @       @               @       @      �?      �?       @�����f�?Щ�-A��?                                SO�o�z�?              �?               @       @       @       @               @      �?      �?       @�`ph>�?2��s4�?                                �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ��?y4��?��&n���?                                ��RO�o�?      �?                                               @       @       @              �?       @�7�B�]�?�r�ة�?      �?                        �'�K=�?      �?       @                       @       @                       @      �?              �?��=���?k��o|��?                      �?        ܥ���.�?      �?       @      �?               @               @       @       @              �?      �?����Z��?5ޫϹ��?      �?      �?      �?        6��9�?      �?       @      �?                                       @                      �?       @1v�z�?w�}��G�?      �?                        v�'�K�?      �?              �?               @       @               @       @                       @�۴���?_m�����?      �?              �?      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @����T�?N@�	�Ǜ?              �?      �?        P�o�z2�?      �?       @      �?               @                               @              �?        �=����?Uin����?      �?                        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        #w\I`ޓ?LE�*AU�?                      �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?        -h#���?fw���?              �?                �'�K=�?      �?              �?                       @               @       @              �?      �?�Gm?C�?�A�Ud�?      �?              �?        ��ۥ���?      �?                       @               @       @       @       @       @      �?       @,���?y�?�JH�w�?      �?                        F���@��?      �?       @      �?                                       @       @                      @���`p�?��q�β?      �?              �?      �?�o�z2~�?      �?       @      �?       @       @                       @       @              �?       @�����?Q�,ߙ��?      �?                        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�d�Q�ϐ?�Z�m�?      �?                      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @^��Z��?_�_�?                      �?        P�o�z2�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�?M��2��?                                ��Vؼ?      �?       @      �?                                                              �?       @HE�����?����?      �?              �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?����[�?��"`�?      �?                        6��9�?      �?       @      �?               @               @       @       @      �?      �?      �?�Dz�rv�?
��r+��?                      �?        Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @����T�?P_]�K��?      �?              �?      �?�]�����?      �?              �?               @       @               @       @      �?      �?      @��_���?3M:z���?      �?      �?      �?        ��ۥ���?              �?                       @       @               @       @              �?        �^<���?�.R����?                                �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        Rp�l?
���*�?              �?                Zas �
�?      �?              �?                               @       @       @              �?       @�Gm?C�?��El�?                                �'�K=�?      �?       @      �?                                                              �?       @84�돗�?oz'��?                      �?      �?�ԓ�ۥ�?      �?       @      �?               @               @               @       @      �?        �H*���?���S��?                                ���V،?      �?       @      �?                                                                      �?�ae��	�? ���U�?                      �?      �?      �?      �?       @               @       @       @       @                       @      �?        ��J��?W���a�?      �?                        $Zas �?      �?                       @               @                       @                      �? .�c�?h\��Qa�?                      �?        (�K=�?      �?       @                       @       @       @       @       @       @      �?        y4��0�?+�����?                              �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @���@��?��5��o�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�Y;���?�]Q�T�?      �?                        P�o�z2�?      �?       @      �?       @       @       @               @              �?                �^<��u�?+1_�0�?      �?      �?                              �?                                                                                       @����e�?���W�g?                      �?      �?H���@��?      �?       @      �?               @                       @       @              �?       @��q%��?=�K���?      �?              �?        �'�K=�?      �?       @      �?       @       @                                              �?       @#���?O�7���?                                [as �
�?      �?              �?       @               @       @                                       @'�F7��?���O���?      �?                        F���@��?      �?       @      �?                                                                       @�Ɉ����?���䓜�?      �?              �?      �?P�o�z2�?      �?       @      �?       @       @       @               @       @       @      �?       @��|�G�?�D�5H��?      �?                      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @n��W�?��H���z?                      �?      �?�D+l$�?      �?                       @                       @               @                        �L�cX��?�M"�?                                ܥ���.�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ��*��?�!g�w�?      �?              �?        p�z2~��?      �?       @      �?                                       @       @      �?      �?      �?��a��?c�����?                      �?      �?p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�bѲ
n�?����U�?              �?                �@�6�?      �?       @      �?               @       @               @       @              �?       @A���Kn�?���!d�?      �?              �?        6���?              �?                                               @       @      �?      �?      �?�{'Y��?r������?                      �?        ��.�d��?      �?       @      �?               @       @               @       @              �?       @)���G��?��v)k��?      �?      �?                p�z2~��?      �?       @      �?               @       @               @       @              �?      �?%��}��?���)�L�?              �?                ,l$Za�?      �?                                       @       @       @       @      �?                ̖p���?�?� ��?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @#w\I`ޓ?�Ր�,%?                                ?���@��?      �?              �?               @                                              �?        =݌S��?v���M��?      �?              �?        p�z2~��?      �?                       @                       @                                      @�����?r!Qn�&�?      �?                        6��9�?      �?       @      �?                                                                       @��C��?=�e�)��?      �?              �?        >�]���?      �?       @      �?               @               @       @       @      �?      �?       @��b�V�?錋�5�?      �?                        6��9�?      �?       @      �?               @                                              �?        �AQ�s��?�����?                              �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @n��W�??3�z�n�?      �?      �?                �@�6�?      �?              �?                                       @                      �?       @�j1v��?h�|��I�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����`�?|�ަ��?                                                      �?                                                                              @����T�?�Ր�,E?                                6��9�?      �?                                                                                      @)g��1�?�B ��7�?      �?              �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @m+�oM�?F��;��?                              �?F���@��?      �?              �?                                                              �?       @�d�Q���?���pjЪ?                      �?        (�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        !�iŽ�?��؞]�?      �?              �?      �?(�K=�?      �?       @               @       @       @       @       @       @       @      �?      �?�
����?&�*&"��?      �?              �?        �
��V�?      �?       @      �?               @       @               @                              �?Y e���?��偯�?      �?      �?                ?���@��?      �?              �?                                                              �?       @�r@��?��q@�?      �?              �?        �]�����?      �?                       @                       @                              �?       @�
����?>�����?      �?      �?      �?        �z2~���?      �?       @      �?                                               @                       @���w���?qbU��?      �?                      �?��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @���C�?]��F��?      �?              �?      �?�D+l$�?      �?                               @       @       @       @       @      �?              �?ï�Dz��?e��³��?              �?                �z2~���?      �?       @      �?                       @               @       @      �?      �?        �
����?;7�6�j�?                              �?ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @8�]�FR�?���s��?                                >�]���?      �?       @      �?               @               @       @       @              �?        AQ�s���?�����?                                F���@��?      �?       @      �?       @                                                      �?      @��<݌�?,)"��N�?      �?      �?      �?        p�z2~��?      �?       @      �?               @       @               @       @              �?       @�N��b�?���@��?                                6��9�?      �?              �?                                               @              �?        !�iŽ�?˾l�o�?                      �?        ���.�d�?      �?              �?       @                       @       @       @      �?      �?      @��!�
�?K��4?�?                      �?      �?��V��?      �?       @      �?       @               @               @       @      �?      �?      @��-�<5�?\?N�0w�?                      �?        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @Y�)L�ْ?G��iiǤ?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                )g��1�?�<�a��?                      �?      �?��RO�o�?      �?       @      �?                                       @                      �?       @y4��0�?=#���?                      �?      �?�RO�o��?              �?                       @                       @       @              �?       @[�՘H�?��܄���?                      �?        ��ۥ���?              �?                               @       @               @       @      �?       @	n��W�?��9���?                      �?         �
���?      �?                               @       @               @       @       @      �?      �?84�돗�?7������?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?                n��W�?��WS�?                      �?        ,l$Za�?      �?       @      �?                                       @       @              �?       @�4�G���?%>U���?      �?                        p�z2~��?      �?                       @       @               @                                        ��V���?�*y� �?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                      @�'�F7�?{����?                                Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?                Y�)L�ْ?ۄ��n��?      �?              �?      �?,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ���@��?�C/`���?                      �?         �
���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����[�?�ųR	�?                                H���@��?      �?                       @                       @       @       @              �?      �?�.M��o�?����(�?                      �?        ��Vؼ?      �?              �?                                               @              �?       @~5&���?8u~�*�?                                �ԓ�ۥ�?      �?                                       @                                      �?      @��e0
8�?�{�C�й?                      �?        �
��V�?      �?       @      �?               @                                              �?      �?��s���?S�Oˊ^�?      �?                        �'�K=�?      �?       @      �?                                               @              �?       @ ʣ��8�?�M��q�?      �?              �?      �?���V؜?      �?                               @       @                                      �?      @z����"�?$K�^˥�?                                6��9�?      �?       @      �?               @                                              �?      �?�����?�T>E��?                      �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @����'t�?��?��?      �?                        $Zas �?      �?              �?       @               @               @       @       @      �?       @
�R,�?VC�#���?                      �?      �?�z2~���?      �?                       @       @               @                      �?      �?      @Alӊ{'�?rq����?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ��w����?4�(���?      �?                      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @9�%��}�?nS�<��s?      �?                        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @-h#���?�|8�?                      �?        �]�����?      �?       @               @                       @       @       @              �?       @��.h�?��u��v�?                      �?      �?��ۥ���?      �?                       @               @               @       @       @              �?�[���?
�LG���?                                ���V؜?      �?              �?                                       @       @              �?       @[ݧ����?��;�0�?              �?                >�]���?      �?       @      �?               @       @       @       @       @      �?      �?       @WH�%���?N�m	��?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?b��1��?W8`�Q�?                                �'�K=�?      �?       @      �?       @       @               @                              �?        d�Q���?o������?                                Zas �
�?      �?              �?               @                               @              �?       @�,u�ئ�?��3��?      �?                        6��9�?              �?                       @               @                                       @۴��I�?��LR�?      �?                         �
���?      �?       @      �?       @       @                                              �?      �?��ds��?>�U,�?              �?      �?        ���V،?      �?                               @                                                      �?��"X~P�?J-?              �?                ?���@��?      �?              �?                                       @                      �?       @���Z�K�?�R��50�?              �?      �?        �RO�o��?              �?                       @                       @       @       @      �?      �?5w\I`��?eu��}U�?      �?              �?      �?SO�o�z�?      �?                       @                       @               @      �?              �?��g{��?�(��D�?      �?              �?      �?��V��?      �?                                       @       @       @       @      �?      �?      @Q�E�*��?JBV�u��?                      �?      �?$Zas �?      �?              �?                       @       @                              �?        +�d�#�?騉�#��?      �?                      �?���V؜?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @���f�´?��w*6�?                                              �?              �?                                       @                               @q
Sb���?C7���|?      �?                        �ԓ�ۥ�?      �?       @      �?                                                              �?        :x��B�?ư�K�S�?      �?                                      �?              �?                                                              �?       @���"X~�?3vA�09x?                                ��Vؼ?              �?               @               @       @       @       @                      @/�Q���?�\�Ȯ?      �?              �?      �?      �?      �?       @      �?       @       @       @               @       @       @      �?        2%fK8O�?�X�]Y�?      �?              �?        �'�K=�?      �?                               @       @                                      �?      @�`ph>�?�t��;�?              �?                SO�o�z�?      �?       @      �?               @       @               @       @              �?        �:Blӊ�?�d�f��?      �?              �?      �?��ۥ���?      �?       @      �?       @                               @       @       @      �?       @��.h#�?��f�r�?      �?                         �
���?              �?                               @       @                                       @۴��I�?3�1�h��?      �?                                      �?       @                                                                      �?      �?፿Po�?8rK��Mm?      �?              �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?      �?                9�%��}�?���'��?      �?                         �
���?      �?                                                                                       @B�]�FR�?o�����?      �?              �?        ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?       @              @]����`�?Is\u��?                      �?        �z2~���?      �?       @      �?       @       @       @       @       @       @      �?              @����C�?�QaT;��?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @^��Z��?�#�`qe�?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?����>u?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�፿Po�?� >�!�[?      �?                        ���V،?      �?                                                                              �?       @<�^!�?����Ղ?      �?                        ���V؜?      �?       @      �?               @       @               @       @              �?        �������?ml(���?                                ��ۥ���?              �?               @       @       @       @               @       @      �?      @}��j1�?6�8���?      �?              �?        {2~�ԓ�?      �?       @      �?                                       @       @              �?        ��vA�?\ݒ��<�?                                F���@��?      �?              �?                                               @              �?       @���Up�?�֏�8̭?                                $Zas �?      �?              �?                       @       @                       @      �?       @*L����?�N+OT��?      �?                         �
���?      �?       @      �?                       @       @                              �?      @�H*���?P�h���?      �?              �?      �?$Zas �?      �?                       @               @       @       @       @      �?              �?M+�d��?`Z��)^�?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?�9�(� ?                                �D+l$�?      �?              �?                               @       @                               @Ͽk�.M�?�|����?      �?              �?      �??���@��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?ò
n�ͭ?��f�<�y?                                ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����`�?w��ٯ�?              �?                �'�K=�?      �?       @                                       @                                      �?jL�*g�?�Q6+Wϵ?                      �?      �?�'�K=�?      �?                       @       @                                                      @�5A .�?�dI�a�?      �?      �?      �?      �?�@�6�?      �?       @      �?               @       @       @       @       @      �?      �?       @WH�%���?ϖ���?      �?                        ��RO�o�?      �?       @                               @       @                                       @H���<�?~�{��?      �?              �?        ��.�d��?      �?              �?       @       @       @       @       @       @       @      �?       @7��+	�?�	��1�?      �?              �?      �?��RO�o�?      �?       @               @       @                               @       @                K��a�?Tt�T�?      �?      �?                ��Vؼ?      �?              �?                                               @              �?       @q
Sb���?��ϫ�?      �?                        Zas �
�?      �?       @                       @       @                       @              �?        5�u�b��?��Rb��?      �?              �?      �?3~�ԓ��?      �?       @               @               @       @               @       @              @����J�?�$�!3�?      �?                        ���V؜?      �?              �?                                               @              �?       @���!���?����ě?                              �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?                �U�����?[��EK�?      �?              �?      �?Zas �
�?      �?       @               @       @               @       @       @                       @ ʣ��8�?O���_�?                                �@�6�?      �?              �?                       @                       @                       @��J��?|\RI�?      �?                        6��9�?              �?                               @               @                      �?       @���vA�?��w���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @�d�Q�ϐ?�9�(� ?      �?              �?        $Zas �?      �?                       @                       @               @      �?      �?      @b/��:�?�1ƛ��?                      �?      �?��V��?      �?       @      �?                                               @                      �?��̱��?w7j#�?              �?      �?        6���?      �?              �?       @       @               @       @       @      �?      �?      �?�����?��4O��?                                �@�6�?              �?                               @               @       @              �?       @{������?52?�?                                ܥ���.�?      �?                       @               @       @                      �?      �?      �?��E�X��?��$i@�?      �?              �?      �?�D+l$�?      �?                       @       @       @       @       @       @       @      �?       @3���?pڊy��?                                ��Vؼ?      �?       @      �?                                       @       @              �?       @&���[�?ߦT����?      �?                        ��.�d��?      �?       @      �?                       @                       @       @      �?      �?[ݧ����?���`���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?       @              @1[�yj�?؄�3��(?              �?                ���.�d�?              �?                       @               @       @                      �?       @z+�oM�?�.Z0�-�?                                H���@��?      �?                                       @       @       @       @       @      �?        �@ʾ���?5U�NY�?      �?                        �ԓ�ۥ�?      �?       @      �?                                                                      �?k� 6\.�?�la�0T�?                                6��9�?      �?                                                               @              �?       @ Q�E�*�? |��?      �?      �?                �z2~���?      �?       @      �?                                                              �?      �?+	�{B��?����?      �?              �?      �?��RO�o�?      �?       @      �?                                                              �?        �ئ�N�?
�M��6�?                      �?      �?�ԓ�ۥ�?      �?       @               @               @       @                       @      �?      �?b/��:�?+��IG�?                      �?        3~�ԓ��?      �?              �?       @                                                      �?        ���I�:�?�����?      �?                      �?�RO�o��?      �?       @               @               @       @       @       @       @      �?       @Ô�-�<�?\���lV�?                      �?      �?,l$Za�?      �?                       @                       @                                        ��s��2�? 4�ߺ�?      �?                        �@�6�?      �?       @      �?                                                                      @���H*�?h�����?              �?      �?        �'�K=�?      �?       @      �?                       @               @       @              �?        ��?y4��?�=�"��?      �?              �?        �
��V�?              �?                               @       @       @       @              �?        �
n���?���V@��?      �?                        �z2~���?      �?       @      �?                               @       @       @              �?      @k1v��?�FQt�?                                ?���@��?              �?                                                                      �?      @b��1��?�!��A�?                                                      �?                                       @                                      @�����T�?���6V?                      �?        �@�6�?      �?       @      �?               @                               @              �?       @,u�ئ�?���-\'�?                      �?        ��ۥ���?              �?                       @       @       @       @       @       @      �?      �?�o��z�?��-d���?                      �?        ���.�d�?      �?       @                               @       @                      �?                �n�)L��?�AYm��?                      �?      �?Zas �
�?      �?       @               @       @                                                       @�^<��u�?;���?                                ���V،?      �?              �?               @                       @                      �?        Ln��4��?�i>��}�?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                       @�%��}�?��߄3�s?                      �?        �V�H�?      �?                               @               @       @               @      �?      �?�ć7�B�?{���<�?                                �K=��?      �?                       @               @       @       @       @      �?      �?        �`�AQ��?F��� �?              �?                ���Vج?              �?                       @                                                       @⛌8j��?�\�k��?      �?              �?              �?      �?       @               @       @       @       @       @       @       @              �?�)����?�}����?      �?              �?      �?F���@��?              �?               @       @       @                               @              @�E�X���?3ۈ�9ݞ?      �?              �?        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                        ��N�ԑ?��.��)m?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                       @�፿Po�?fN
u�w*?              �?                ���Vج?      �?              �?                       @               @                      �?      @<��u�4�?(�Y�p�?                                6��9�?              �?                       @                               @              �?       @�#�d�Q�?�y�<�k�?      �?      �?                                      �?                       @       @                       @              �?       @j?C؋��?�i��(g?                      �?      �?3~�ԓ��?      �?                       @       @               @                                        �o��z�?/3�C�?      �?      �?                $Zas �?      �?              �?                                                                      �?�Z�<��?R���=�?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�'�F7�?�	� �?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ���Z��?��2���?      �?                        ��Vؼ?      �?              �?                                               @              �?       @�:]���?��-����?      �?                        �z2~���?      �?       @      �?                                       @                      �?       @#���?o��Ș��?      �?                        ���Vج?      �?              �?                                       @                      �?       @r�g�L��?(�Y�p�?                                �@�6�?      �?              �?                                                                      �?@y4���?�a_x��?      �?              �?        �'�K=�?      �?       @      �?                       @       @       @       @       @               @_�ti���?ߡ]���?                      �?      �?���.�d�?      �?       @      �?       @       @               @       @       @       @                2%fK8O�?�������?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        E�(Ţe�?��w���?                                ���V؜?              �?                                               @                              �?�����?��o�N�?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @                #w\I`ޓ?�� ��?      �?              �?      �? �
���?      �?              �?                                               @      �?                L���S�?������?                                �@�6�?      �?                                       @       @               @      �?              �?@�MF��?_�~��
�?      �?              �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                       @F��1��?��UR�g�?              �?      �?      �?�o�z2~�?      �?       @      �?               @       @                       @              �?      �?�4�G���?\c@W(�?              �?                              �?              �?                                                              �?       @돗�(��?;ⴴc�x?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?                      �?��N�ԑ?F�eP�A�?      �?                        ��Vؼ?      �?              �?                       @               @       @              �?       @z����"�?�?.��k�?                      �?        v�'�K�?      �?       @      �?       @       @               @                      �?               @�F��?�T�2��?                                H���@��?      �?       @               @       @       @       @       @                      �?        &`��"�?���h��?      �?                        �ԓ�ۥ�?      �?       @               @                                                              @��s��2�?FF�=?�?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�፿Po�?������?      �?      �?                �6��?      �?       @      �?                                       @       @                       @&���[�?�ȅ���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @����[�? �<$3?                                �z2~���?      �?              �?                                               @                        V����?ضm۶m�?                                (�K=�?      �?       @               @       @       @               @       @       @              @��a�(�?Ó���?      �?                      �?              �?              �?                                                                        ����e�?M�$&�x?                                H���@��?              �?                               @               @       @              �?       @�rv��?7[�:��?                              �?              �?              �?                                       @       @              �?       @�G�Ɉ��?����;��?              �?                �@�6�?      �?       @      �?                                       @       @              �?       @��s��2�?!!����?                                              �?              �?                                                              �?       @cX�~k��?EF�=?x?                                �@�6�?      �?       @      �?                               @       @                               @�
����?V�� ��?      �?      �?                6��9�?      �?              �?       @                                       @              �?       @�Ήo��?�����?      �?              �?        3~�ԓ��?      �?       @               @                       @       @              �?      �?      �?�<�^�?jQV�?                              �??���@��?      �?       @      �?               @       @                                                
Sb����?�C�`���?                      �?        ��V��?      �?              �?       @               @       @       @       @      �?      �?       @Wc"=P9�?O����?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?nC��x�?D�%�>�v?                                �z2~���?      �?       @      �?                                       @       @              �?       @����?d�^Gh'�?                      �?        F���@��?      �?              �?                                                              �?        �c9�?X�k��?      �?      �?                ���V،?      �?       @      �?                                                              �?      @�ht3N�?A:���?      �?              �?      �?P�o�z2�?      �?              �?               @       @       @       @       @      �?              �?�b�V��?\OD�6��?      �?              �?      �?              �?              �?                                               @                       @M+�d��?��!�|?      �?      �?      �?              �?      �?       @                       @       @       @       @               @              �?�0@�b��?�R}R��?                      �?        �@�6�?      �?       @                                                                               @���7q�?T�C-y�?      �?                      �?,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?       @                �%��}�?%�����?              �?                              �?              �?                                       @       @              �?       @}�mu��?�>�5��?      �?                      �?�]�����?              �?               @       @       @                                      �?       @��>�MF�?�E����?                      �?      �?SO�o�z�?      �?       @       @      �?      �?      �?      �?      �?      �?       @               @M:'>��?�/0�h�?      �?      �?      �?              �?              �?               @       @       @       @       @       @       @      �?      �?��Ͽk�?nd��y�?      �?                        ��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�rv��?�Im�)�?      �?              �?        �'�K=�?      �?              �?                       @                                      �?      �?���H*�?`
���?                                              �?              �?                       @                                                84�돗�?,L�
��y?      �?              �?        �ԓ�ۥ�?      �?       @                       @                                                      �?JS}䛌�?�H�0�?      �?              �?      �?(�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?n��W�?�h7O��?                                ��Vؼ?      �?              �?       @                                                      �?       @̖p���?�Z�]�?      �?              �?        p�z2~��?      �?       @      �?               @       @                                      �?        ^<��u��?������?                      �?      �?              �?              �?                                                              �?      @%�yO�0�?#��=�w?      �?              �?      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�m��W�?60��H�?                                6��9�?      �?       @      �?                               @       @       @              �?       @P9��_��?ʱ8Ĵ�?              �?                {2~�ԓ�?      �?              �?                                       @       @              �?       @^!ї�V�?V��T���?                      �?        �RO�o��?              �?               @       @               @                       @                �i����?�ek}��?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?       @��(��|�?�h����?                      �?        �6��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�����`�?z� �P��?                              �?���V،?      �?       @      �?       @                                                              �?��r�9��?�g�F�?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @E�(Ţe�?�}xK�Θ?      �?                        �D+l$�?      �?       @      �?       @       @       @       @                              �?      �?���`p�?�"R9��?      �?              �?      �?>�]���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �^W-��? U&�o�?                      �?        �K=��?      �?       @      �?       @               @       @       @       @      �?      �?       @�1����?rPh��?                      �?        ��ۥ���?      �?       @      �?       @               @               @       @      �?      �?      �?�����U�?��=�M�?                      �?      �?�D+l$�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @\��r�?�d	ŽĶ?      �?      �?      �?              �?      �?       @      �?               @       @       @       @       @       @      �?        Ň7�B��?+���A��?                      �?      �?�z2~���?      �?       @      �?               @       @                                      �?       @�s��2�?���ч�?                                �z2~���?              �?               @                       @                      �?      �?      @��<݌�?lj1jŝ�?                      �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @M:'>��?K��捷�?                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @                Y�)L�ْ?Zxv�L�?                      �?      �?H���@��?              �?               @                       @                      �?      �?      �?�R,Z�?�ųR	�?                      �?      �?�@�6�?      �?                                                       @                               @؋�ߵN�?w\�.}ޣ?              �?                �'�K=�?      �?       @      �?                               @       @       @              �?      �?w\I`��?]Ĕ��H�?      �?              �?        �
��V�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ��+$��?[ł���?      �?                        p�z2~��?      �?       @      �?               @       @               @       @      �?      �?       @o��T�?z�o���?      �?                        �]�����?      �?       @      �?               @                                              �?       @��+$��?;:����?      �?      �?      �?                      �?       @      �?                                       @       @              �?       @{]�;x�?|qU!�?      �?              �?      �?6��9�?              �?               @               @       @                      �?      �?       @h�����?�W~�@�?      �?              �?      �?���@��?      �?       @      �?               @               @       @       @                       @��-�<5�?�y���?      �?              �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              @-h#���?#LT�nX�?      �?                        �ԓ�ۥ�?      �?       @      �?               @       @       @       @               @      �?      �?[�yjH�?-C�����?      �?                        ?���@��?      �?       @                                                                              �?UUUUUU�?J������?      �?                        ��Vؼ?      �?       @      �?       @                                                      �?       @�b��!�?1��C,��?                      �?        H���@��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      @��dsǵ?k���>�?                                �@�6�?      �?              �?                                                                        ��w����?9>��
�?      �?      �?      �?        Zas �
�?      �?              �?               @                                              �?      �?j�����?%
��  �?      �?                        6���?      �?               @      �?      �?      �?      �?      �?      �?       @              @ś�8j��?]<+����?                                �D+l$�?      �?              �?                       @               @       @       @               @'t J��?/��JX��?                      �?        �]�����?      �?              �?                                                              �?       @o�Wc"=�?%u�m��?      �?                        ���V؜?      �?                       @               @               @       @              �?       @��4�u��?Y�H#�?                                �z2~���?      �?       @      �?                                               @              �?       @&�1�L��?���?.��?                                [as �
�?      �?       @      �?       @               @                                      �?      �?�iŽ�,�?�b�l^)�?                                �@�6�?      �?       @                               @       @               @      �?      �?       @���&�?ߞ����?      �?              �?      �?6��9�?      �?       @      �?                       @       @       @       @                       @{B���?D4�\s�?                                ��Vؼ?      �?                                               @       @                      �?        ��¯�D�?}�"�4�?                                �'�K=�?      �?       @      �?               @               @               @      �?               @c9�W�?QyŸ �?                      �?        3~�ԓ��?      �?              �?               @                               @                        ��Kn���?|!.�x��?      �?      �?                ��Vؼ?      �?       @      �?                                               @              �?      �?a�:�?�o�N�?                      �?      �?�ԓ�ۥ�?      �?       @               @       @                                              �?      �?H���<�?P�.?�H�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      �?E�(Ţe�? ��??                      �?      �?v�'�K�?      �?                       @       @               @                       @      �?      �?��	�p�?v�B.�?      �?              �?      �?�V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @Y�)L�ْ?��ٯ�?      �?      �?      �?        6��9�?      �?       @      �?                       @                       @              �?       @�hY7��?`Ugw't�?                                [as �
�?      �?       @      �?                               @                              �?      �?��*��?��c�?      �?                        6��9�?      �?       @      �?       @                               @                      �?       @F�*�A6�?*W�Ub��?                                3~�ԓ��?      �?       @      �?               @       @       @       @       @              �?      �?S��*�?�/v.$��?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?E�(Ţe�?��ټ�?                                6��9�?              �?                                       @                       @      �?      @$X~PT�?�wɦ���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                       @8�]�FR�?����d!?                                ?���@��?      �?       @      �?               @               @               @              �?       @����?����I�?      �?                        �]�����?              �?                               @       @       @       @       @                ƽ�,u��?�!����?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?�W�ħJb?      �?                      �?�'�K=�?              �?                                                                              @�6��w�?7�r5�?                      �?        �V�H�?      �?                       @       @               @               @      �?              @D)-��?M�O,��?      �?                        ,l$Za�?      �?       @      �?       @       @       @               @       @              �?       @z'Y���?8S]f��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?�^/��"?                                6��9�?      �?       @      �?                                               @                       @�WH�%��?������?      �?              �?      �?�'�K=�?              �?               @       @       @       @               @      �?      �?      �?c9��?D�C���?                      �?      �?�ԓ�ۥ�?      �?       @               @               @       @       @                               @*g��1�?	�#;���?              �?                Zas �
�?      �?       @      �?                                       @       @              �?       @~�ɣ���?�A%O�?                                ���V،?      �?                                       @       @       @       @                       @m$���?�V�uǐ?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?���i�A�?      �?              �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @m+�oM�?ѣw�@G�?                              �?���V،?      �?       @      �?                                       @       @              �?        ���.�?�p���?      �?                                      �?                       @                                                              @~5&��?Tab:Ӭn?                      �?      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?                      @�'�F7�?0�P�_�?                                �6��?      �?       @               @       @       @               @       @      �?                �W���?�j��g�?      �?              �?      �?�ԓ�ۥ�?              �?                       @       @               @              �?              �?8ֳv&��?����q�?      �?              �?        $Zas �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����'t�?�y�G��?      �?                        6��9�?      �?       @                               @       @                                       @!s�g�L�?<����?      �?                        H���@��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�d�Q�ϐ?bRD*��?      �?      �?      �?      �?�ԓ�ۥ�?      �?                               @               @       @       @              �?       @�c=kg�?�x�U&�?                                �'�K=�?      �?       @      �?       @                       @       @       @              �?        ?|]��?q��xy�?                      �?      �?      �?      �?                       @       @       @               @               @      �?      �?�r@��?�v�-Io�?      �?              �?      �?��ۥ���?      �?       @      �?               @                       @       @      �?                ���?y4�?Gr���2�?      �?                        Zas �
�?      �?       @                       @                                                       @��W��?/M��M�?                      �?      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?                        m+�oM�?{����?                      �?      �?���V،?      �?              �?                                                                       @�V�ߚ�? ���U�?              �?      �?        ��V��?      �?       @      �?               @       @               @       @              �?        Tb�����?�}�J�?      �?              �?      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��C��?"�0��?      �?                                      �?                                                       @       @              �?      @8j��^�?�� ��t?                      �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�'�F7�?��O���?                              �?              �?              �?                                       @                      �?       @d��ht�?����z�|?      �?      �?      �?        $Zas �?      �?       @      �?                                       @       @              �?       @�0%fK�?�f�o���?                                              �?              �?                                                                       @cX�~k��?EF�=?x?      �?                        $Zas �?      �?       @      �?                                       @                      �?       @UUUUUU�?����mW�?      �?      �?      �?        �o�z2~�?      �?       @      �?       @       @       @                                      �?       @R��'��?���:��?      �?                        F���@��?      �?       @      �?                                               @              �?      @��`�AQ�?q<�8�>�?      �?              �?        H���@��?      �?              �?                       @       @       @       @      �?      �?      �?����?�ӯ��?      �?                      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�፿Po�?����^�?                      �?      �?�'�K=�?      �?                       @                               @       @      �?      �?        cX�~k��?)�$���?                                              �?                       @       @                                              �?       @]!ї�V�?�C��q?      �?                        3~�ԓ��?      �?       @               @       @       @       @                      �?                ���'t�?��ROg9�?                      �?      �?��V��?      �?       @      �?       @               @               @       @       @      �?      �?��0%f�?p������?              �?                �@�6�?      �?       @      �?                                               @              �?      �?y4��0�?$�jg�;�?                      �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�]�FR�?�}U�ݝ�?      �?                                      �?                       @                                                      �?      @���Z�K�?h�Zlnl?      �?                                      �?              �?       @                                       @              �?      @l	�Y �?w�\�?      �?              �?        �@�6�?      �?       @      �?               @       @       @       @       @              �?       @�f���?�v�.��?                                ���V؜?      �?              �?                               @               @                       @��H*��?�K��F�?      �?      �?      �?        ���Vج?      �?       @      �?                       @                                      �?        ȕ�=��?�M%��5�?      �?      �?      �?      �?              �?                                               @                              �?      �?!�iŽ�?|��h��l?                                �@�6�?      �?              �?               @               @       @       @              �?        9�)1[��?����z��?      �?                        �'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @�{B���?U�eP�A�?      �?                                      �?       @                       @                                                       @����?�V�u�p?                      �?        >�]���?      �?       @      �?               @                       @       @      �?      �?       @�C��x�?�KnJE�?      �?              �?        ���Vج?      �?       @      �?       @                                       @              �?       @��Y;��?ـ���M�?                                              �?                                                                                      @��}�ɣ�?��f�<�i?      �?                        ���V؜?              �?                       @               @                              �?      @"��~���?����>�?      �?              �?                      �?              �?                                                                       @�¯�Dz�?Ӧ<$3x?              �?      �?        ���Vج?      �?              �?                                                              �?       @�vAIE�?�)�M�?                      �?      �?��RO�o�?      �?              �?                                               @              �?        m$���?�����?      �?              �?      �?SO�o�z�?              �?               @               @       @       @               @              �?�G��q
�?�iy��?                                $Zas �?      �?              �?       @               @       @       @              �?      �?       @X~PT��?���=/"�?                                              �?               @      �?      �?      �?      �?      �?      �?                      @F��1��?��ֺ�?                                �z2~���?      �?                                       @                                              �?�b��!�?�����b�?                                �RO�o��?      �?               @      �?      �?      �?      �?      �?      �?       @                m+�oM�?�L�(�b�?      �?                      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�X����?+�^�?                                !�
���?              �?                       @       @               @       @      �?      �?      �?�0%fK�?��^}�?      �?      �?              �?              �?                                       @                                      �?      @��"X~P�?�Ŏ���m?                                $Zas �?      �?              �?       @               @               @                      �?        ��%���?ȼ7�!\�?                      �?        �RO�o��?      �?       @      �?               @       @               @       @              �?       @�g{���?ߎ�%Κ�?                                6���?      �?       @               @       @       @       @                      �?      �?      �?�/�����?���׍��?      �?      �?      �?        �V�H�?      �?       @      �?                       @               @       @              �?       @��l	��?�!L�q��?                      �?              �?      �?       @      �?               @                       @       @       @      �?      �?�n�)L�?�0�-L�?      �?              �?              �?      �?       @      �?       @       @       @                       @       @      �?       @9�)1[��?W'��]V�?                      �?        F���@��?      �?       @      �?               @       @               @                               @=���&�?NZ[��?                                              �?                                                       @                      �?      �?jL�*g�?�ᙁ(q?      �?                        ���Vج?      �?                               @               @               @              �?        �U:'�?I��W���?      �?      �?      �?        !�
���?      �?       @      �?       @               @               @                      �?        ����C�?0��`Qy�?                                ��RO�o�?      �?                               @       @       @       @       @      �?              @ݧ����?V�.�m�?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @              @�L�5A �?�qpTV��?                      �?        �@�6�?      �?                                                                              �?       @�bѲ
n�?v���w�?      �?                        ���V،?      �?                                               @       @       @                       @p�l�?XIW�؊?                                �z2~���?      �?                                                                                        �vAIE�?���qٮ?                                	��V��?      �?       @       @      �?      �?      �?      �?      �?      �?                      @�r@��? ���?      �?                        P�o�z2�?      �?       @               @       @       @                       @      �?      �?      �?�X���??^��|z�?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @8�]�FR�?����ě?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �X����?)ɀM�y�?      �?                        ܥ���.�?      �?                               @       @       @       @       @       @              �?��䶺O�?=�z��?              �?      �?        6��9�?      �?       @      �?                                                              �?       @��x��?�>�? �?                                e�v�'��?      �?       @      �?       @               @               @       @      �?      �?        e����I�?TKy����?      �?                      �?$Zas �?      �?               @      �?      �?      �?      �?      �?      �?              �?       @�፿Po�?��C��?              �?      �?        e�v�'��?      �?       @      �?               @                       @       @      �?      �?      �?���?�r3>p��?      �?                        ?���@��?      �?                                       @       @       @       @              �?       @�u�b���?`Hqm���?                      �?      �?      �?              �?               @       @       @       @               @       @              �?;�^!��?�o-��?      �?                        �@�6�?      �?              �?       @                                                      �?       @84�돗�?����`ն?                                F���@��?      �?                       @       @               @       @       @              �?       @ph>�/�?a���YP�?                      �?      �?6��9�?      �?       @      �?                                       @       @              �?       @Ž�,u��?��06V�?      �?              �?      �?�o�z2~�?      �?               @      �?      �?      �?      �?      �?      �?      �?                8�]�FR�?�����?              �?      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?�Q���\�?o��p�~�?      �?                        ��RO�o�?      �?       @      �?                               @       @                      �?       @��7q��?�}]� �?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @                -h#���?7�����?      �?              �?      �?�D+l$�?      �?       @               @       @       @       @                                       @�|�Gm�?͡��D�?                                ,l$Za�?      �?       @      �?               @       @                                      �?        y4��0�?��Bc�?      �?                        p�z2~��?      �?                       @       @       @       @       @       @      �?      �?        ?C؋���?*	�a}m�?      �?                        ��ۥ���?              �?               @       @       @       @       @               @                g{����?[�]��?      �?      �?                �
��V�?              �?                               @               @       @      �?      �?        yO�0@�?��>�?              �?                p�z2~��?      �?       @      �?               @               @       @                      �?       @����'t�?h��%e��?      �?                        ���.�d�?      �?              �?       @       @                       @       @      �?      �?      �?��'t �?�?|��P�?      �?              �?      �?      �?      �?                       @               @       @       @       @       @      �?       @�:]���?a��Rr�?      �?              �?      �?              �?              �?                                                              �?      @�r@��?�+{Hʁx?                      �?        ���V،?      �?                                                                              �?       @�{'Y��?5&�oĀ?                                v�'�K�?              �?               @               @       @       @       @       @      �?        z�D_r�?j�!���?      �?              �?      �?�D+l$�?      �?       @      �?                                       @                               @b�(Ţe�?\���e�?      �?                                      �?       @                                                                      �?       @��"X~P�?�Ŏ���m?      �?                        ���V،?      �?       @      �?                                               @              �?       @�6��w��?f^�T�?              �?                ��ۥ���?      �?       @      �?                                                              �?        �ae��	�?×Tin��?                      �?        �z2~���?      �?                       @               @       @               @      �?      �?        ����`�?͖���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @#w\I`ޓ?�Ր�,%?                                F���@��?      �?              �?                       @                                      �?       @_W-��?F�3�?      �?              �?        ,l$Za�?      �?                               @       @       @       @              �?      �?       @Y�ڙ���?:������?                      �?      �?�K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�j1v�?��)CL��?      �?                        6��9�?      �?              �?               @                                              �?      �?��Po��?�5��@��?      �?              �?      �?��.�d��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�r@��?�%:g��?      �?                        ���Vج?      �?                                               @                              �?       @��̱���?��wh�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?      @n��W�?_�]Q�Tc?      �?                        �o�z2~�?      �?       @      �?                       @               @       @      �?      �?       @��C���?�T���?      �?                        6���?      �?              �?       @       @                       @       @      �?                9�)1[��?_��#C�?      �?                                      �?       @      �?                                                              �?       @���H*�?sn:Oo�z?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?       @       @       @       @       @       @       @      �?        �L�cX��?�G
Z�<�?      �?                                      �?                                                                                      @?y4���?_�<$3h?      �?              �?      �?��RO�o�?      �?       @      �?               @               @                              �?      �?��`�AQ�?��
����?                                �RO�o��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @)g��1�?>S�G���?                      �?      �?      �?      �?       @               @               @       @                       @                ���J��?J։���?              �?      �?        ܥ���.�?      �?                               @                               @      �?      �?        �p����?�WlϮv�?              �?      �?        �ԓ�ۥ�?      �?       @      �?       @       @               @       @                      �?        ����e0�?`O�l���?      �?              �?      �?�D+l$�?      �?       @      �?       @       @                       @                      �?       @�FR,?�?%���R��?                      �?        p�z2~��?      �?       @      �?       @       @       @               @                      �?       @ /�Q���?��Ta��?              �?      �?        (�K=�?      �?       @      �?               @               @       @       @       @      �?        z�D_r�?z|�.��?      �?      �?                �'�K=�?      �?              �?                                                              �?       @K��a�?���6�?      �?                         �
���?      �?                                               @                                        ���w��?Ç^�h��?      �?                        e�v�'��?      �?              �?       @       @               @       @       @      �?      �?      �?��Ͽ�?"�8���?              �?                �@�6�?      �?       @      �?       @       @       @               @       @              �?       @e� �;�?��:?�?                                F���@��?      �?       @               @               @               @       @              �?       @?^��C�?���ټ?                      �?        (�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                -h#���?h�8�]�?                      �?      �?[as �
�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�%��}�?tI���?      �?              �?      �?!�
���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�%��}�?��{K��?      �?                        H���@��?              �?                               @                                      �?        FaJ̖p�?�,�(e/�?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?              �?      @��1�~? �<$3�>                                              �?       @                                                                      �?      @9�WH�?(���m?                      �?      �?��ۥ���?      �?       @               @       @       @       @                       @              @�/�����?8�Hd9�?                                e�v�'��?      �?       @      �?                       @       @               @       @      �?        {]�;x�?��Qt��?              �?      �?        6���?      �?       @      �?                               @       @       @              �?        GR,?(�?:�
ƈ)�?              �?      �?        F���@��?      �?              �?                                                              �?       @'#��~��?�����?      �?              �?      �?���Vج?      �?              �?       @               @                       @              �?      @����?j��g��?                                $Zas �?              �?                               @               @       @              �?       @ئ�N��?�K�grn�?              �?                3~�ԓ��?      �?              �?                                               @              �?       @�?^���?�����?      �?              �?        ���V؜?              �?                       @                                                      �?��Ͽk�?7�3��݁?      �?                        e�v�'��?      �?       @      �?       @       @               @       @       @       @      �?      �?!�iŽ��?n��r�3�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                        �'�F7�?.��2��?              �?                �'�K=�?      �?              �?                       @               @       @              �?       @��U����?1#E�?      �?              �?                      �?                                                                                      �?f��	��?]v�{h?              �?                �'�K=�?      �?       @      �?                                                              �?      @�@ʾ���?�3���?                      �?        	��V��?      �?       @                       @                       @       @              �?        /M��o2�?�����A�?                                ���Vج?              �?                       @                       @       @              �?      �?�������?��ؖ�?      �?      �?      �?      �?�]�����?      �?       @      �?               @       @       @       @       @              �?        F��s�?N��l�=�?                                              �?              �?               @                                                       @G��q
S�?�j)��z?                                F���@��?      �?              �?                                       @                      �?      @EDDDDD�?�AX��ֽ?      �?      �?                �z2~���?      �?       @      �?                                       @       @              �?        1[�yj�?�<�z��?                                �z2~���?      �?              �?       @                               @              �?      �?      �?Ͽk�.M�?��\E�]�?      �?      �?                ���Vج?      �?              �?                                                              �?      @��j1v��?����ؤ?      �?                        F���@��?      �?                                               @                              �?      @�Po���?݇VE�|�?                      �?        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              @���C�?���)*�?      �?                        ���V؜?      �?                       @                                                      �?      @��"X~P�?�����Ȑ?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?b��1��?�I�L}�?                      �?        ��Vؼ?              �?                               @               @       @              �?       @�I�:Bl�?C�b*��?                      �?         �
���?      �?                               @               @       @       @              �?       @\��r�?L9�3��?      �?                        ���V؜?      �?              �?                       @                                      �?      �?�Ɉ����?ީ�]@�?      �?                        p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @              @nC��x�?{Ν�6��?              �?      �?        �'�K=�?      �?       @      �?                                               @              �?       @G�mZq��?v6����?                      �?      �?Zas �
�?      �?       @      �?       @       @       @                       @      �?      �?      �?��S�@�?��fڭ'�?      �?      �?      �?      �?��ۥ���?      �?       @                       @       @       @               @      �?      �?        �%��f�?�����?                      �?        �V�H�?      �?       @      �?               @       @       @       @       @       @      �?      �?���<��?�����?      �?              �?        	��V��?      �?              �?                                                              �?        �V�ߚ�?l�P�~��?      �?                        ���Vج?      �?                                       @               @       @      �?      �?      @�¯�Dz�?���j�?                      �?      �?��Vؼ?      �?                               @               @       @              �?      �?      @�U:'�?��d���?                      �?        �@�6�?      �?       @      �?               @                       @       @              �?       @�������?[& ���?      �?              �?        ���.�d�?      �?       @      �?       @       @       @                              �?                [ݧ����?R�����?                                ��.�d��?      �?       @      �?       @       @               @       @       @      �?      �?      �?�1����?��a���?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?B6w\I`�?˽��?      �?                      �?���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      �?E�(Ţe�?x c[�c�?                      �?      �?�o�z2~�?      �?       @      �?               @       @       @       @       @      �?      �?       @����w�?�s,� 1�?      �?                        �ԓ�ۥ�?      �?                                       @       @                                      �?��J�ć�?�ʇ����?      �?                        �@�6�?      �?       @      �?                                                              �?       @�ae��	�?�h�XO��?              �?      �?        �K=��?      �?                                       @       @       @              �?                �ć7�B�?Q���H��?      �?              �?        ���@��?      �?       @      �?                               @       @       @      �?               @	{�����?��!D:��?      �?                        v�'�K�?              �?                                       @                      �?              �?�U�����?8b����?                                              �?                                                                                       @<�^!�?M�̡��h?                                {2~�ԓ�?      �?       @      �?               @       @               @                      �?        �o2���?�.�%U��?              �?      �?      �?�D+l$�?      �?       @      �?                       @                       @              �?      �?��Dz�r�?K?fS��?      �?                      �?6��9�?      �?                       @       @               @                       @              �?�X����?���K��?              �?      �?                      �?              �?                                                              �?       @���U�?�^��w?      �?              �?        �K=��?      �?       @      �?       @       @       @               @       @      �?              �?Ͽk�.�?п7R��?      �?                        �D+l$�?      �?                                       @                       @      �?      �?        z�D_r�?.�b���?      �?                                      �?                                                                              �?      @�?���}p�h?      �?              �?      �?���V،?      �?               @      �?      �?      �?      �?      �?      �?      �?              @m+�oM�?��)*`?                                �RO�o��?              �?               @               @               @       @       @               @�����?��8%r��?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?              �?      @]����`�?xjD",�?      �?              �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�r@��?�4��
h�?      �?              �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @���6�?)��!D�?      �?              �?        {2~�ԓ�?      �?                               @                                              �?      @��"X~P�?O�BŊ �?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����'t�?nWʜKa�?                                ���Vج?      �?              �?                               @               @              �?      �?��3i�a�?]��*T�?      �?                        ��Vؼ?              �?                                               @       @              �?       @�'t J�?>;�:�?      �?                        �'�K=�?              �?               @                                                              @��>�MF�?�� �Z�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @����'t�?�Z �2c�?              �?                ��RO�o�?      �?       @      �?               @       @                                      �?        �WH�%��?U?��?      �?      �?      �?        F���@��?              �?               @                                                                ��Ͽk�?G�0��ӗ?      �?                        ���.�d�?      �?       @      �?                       @       @       @       @      �?      �?      �?�X����?.)�$._�?              �?                �'�K=�?      �?       @               @       @                                              �?        ��l	��?bBN���?                                ��V��?      �?       @      �?       @       @               @                      �?      �?       @t3NaJ��?r�3A2��?      �?                        ,l$Za�?              �?                       @       @               @       @      �?      �?      @g{����?˲Ņgg�?              �?      �?                      �?              �?               @                                              �?      @m$���?�;���9{?      �?              �?      �?              �?              �?                                                              �?      @X-�r�?�3�
'x?                      �?      �?�]�����?      �?       @      �?                                                              �?        G��q
S�?2���?      �?                        ��RO�o�?      �?       @                       @       @       @               @       @      �?        Q�E�*��?(�ԝ��?      �?              �?      �?P�o�z2�?      �?       @                       @       @       @               @      �?      �?        G��q
S�?��) �z�?                      �?      �?      �?              �?               @       @       @       @       @       @       @                �J�ć7�?&���R��?      �?                         �
���?      �?              �?                       @       @       @       @              �?       @�������?��8-��?                                �D+l$�?      �?                       @       @       @       @       @       @      �?                ��>|]�?C���r��?              �?                ��Vؼ?      �?              �?                                       @                      �?       @B�/����?{�� ��?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?              �?      @E�(Ţe�? ��??                                �z2~���?      �?              �?                       @               @       @              �?       @4�돗��?�֟��Ѿ?      �?              �?      �?$Zas �?      �?       @      �?               @               @       @                              @fK8O��?�!����?                      �?              �?      �?       @      �?               @       @       @       @       @      �?      �?       @/�Q����?��Ss��?      �?              �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�፿Po�?<������?                              �?F���@��?      �?       @      �?               @       @               @       @      �?      �?      �?q���Y�?pI����?      �?              �?      �?�ԓ�ۥ�?      �?              �?               @               @       @              �?      �?       @+�oM��?*G٬\=�?      �?              �?      �?�]�����?      �?       @      �?                       @               @                      �?       @��Dz�r�?w�!���?                      �?      �?(�K=�?      �?       @               @       @       @       @       @               @               @�AQ�s��?Vp�`��?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                        ]����`t?���sO<p?      �?              �?              �?      �?       @      �?       @       @               @       @       @       @      �?      �?ۙ�ǰ2�?��!��?                                ��.�d��?              �?               @       @       @               @       @       @      �?        ����?$V�)M�?      �?              �?        3~�ԓ��?      �?       @      �?                       @                                      �?       @��䶺O�?��>c���?              �?                	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����'t�?��$�k�?                      �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @                8�B�]��?��4Z�?                      �?        3~�ԓ��?      �?       @               @       @                       @       @      �?      �?      �?�j1v��?�c�����?              �?                �@�6�?      �?              �?                       @                                               @�u�b���?5/�CZ��?                      �?              �?              �?                       @       @               @       @       @      �?       @�
����?�G5����?                      �?      �?6���?      �?       @      �?       @       @                               @              �?        �o2���?�iF� �?              �?      �?      �?ܥ���.�?      �?              �?       @               @       @       @       @              �?       @�Dz�rv�?|8����?                                �'�K=�?      �?                                                                                      @�r@��?��C��?              �?                �D+l$�?      �?       @      �?       @       @       @                                              �?����c�?v��;�?      �?              �?      �?6���?      �?                               @               @       @       @      �?      �?      �?""""""�?UZC<���?              �?                �V�H�?      �?              �?               @                       @       @      �?              �?Ž�,u��?�g�pD�?      �?              �?      �?�D+l$�?              �?               @               @                              �?              @ ���?2�w����?      �?      �?                6��9�?              �?                       @       @                                               @�፿Po�? X�5%�?              �?      �?        �@�6�?      �?       @      �?                                               @              �?       @����?湫[r�?      �?              �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @nC��x�?�)�-��?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      �?n��W�?��T#�?                                �@�6�?      �?              �?               @       @                       @              �?       @�^!ї��?����<�?      �?                      �?              �?                               @                                              �?       @���'�?Ѯ^� fm?      �?              �?      �?v�'�K�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�k�.M��?�0�"ml�?                                p�z2~��?      �?              �?       @               @       @       @       @      �?      �?       @��-�<5�?z�̹f�?                                �o�z2~�?              �?                       @       @                       @       @      �?      �?� �;�$�?����*)�?      �?      �?                ��Vؼ?      �?       @      �?                                               @              �?       @H*��E�?ܘ��-�?                      �?      �?�ԓ�ۥ�?              �?                       @       @               @       @       @      �?      �?䶺O_�?�`QyŸ�?      �?              �?        �z2~���?      �?       @      �?       @       @       @               @                      �?       @����?5�e�?      �?              �?      �?      �?              �?               @       @       @       @               @       @      �?      �?#��~���? ��e���?                      �?        >�]���?      �?       @      �?                       @       @       @       @       @                ���I{�?�k��a$�?      �?              �?      �?�RO�o��?      �?                       @       @               @       @       @              �?      �?����[�?B&{�&�?      �?              �?      �?�K=��?              �?                               @       @       @                      �?       @��j1v��?h��A��?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?޵�8�o?                                p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�፿Po�?�dI�a�?      �?              �?      �?�RO�o��?      �?                               @               @       @       @       @                �ڙ�ǰ�?�cFۣ��?                              �?F���@��?      �?       @               @       @       @       @       @       @       @              �?�����?�q����?                                6���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�bѲ
n�?rA=��(�?                                �@�6�?      �?       @                                                       @              �?      @�p����?p�/
b7�?                                �'�K=�?      �?                       @               @       @                                       @�p����?���O��?      �?              �?      �?�@�6�?      �?       @      �?                       @       @       @       @      �?      �?       @�+$����?����>��?      �?                      �?�]�����?      �?              �?               @       @               @                      �?       @��%���?��KI�?      �?              �?      �?[as �
�?      �?       @               @       @               @               @      �?      �?        ��~5&�?^B��,�?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                        �����`�?X�gI<�?              �?                ���V،?      �?       @      �?                       @                       @              �?       @��q
Sb�?�4R���?                                !�
���?      �?       @      �?       @       @       @               @       @      �?                �����f�?���!g��?                                ?���@��?              �?               @                                                      �?      @=Q�s�û?ql�����?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @�፿Po�?���A��?                                F���@��?      �?       @      �?       @                                                      �?      �?M+�d��?�j$6ڽ?                                ���V؜?      �?       @      �?                                                              �?       @S,ZV��?V/X��?              �?                �V�H�?      �?       @      �?       @       @       @               @       @      �?      �?       @�d�#�6�? �d��?                      �?      �?      �?      �?                       @       @       @       @       @       @       @                 J�hY�?���.��?              �?                              �?       @      �?                                                              �?       @�J���?���V/z?      �?              �?        �ԓ�ۥ�?      �?       @      �?                               @       @                      �?      �?�V�;�R�?k�?Y��?                      �?        �K=��?      �?       @                       @       @       @       @       @       @                ��̱��?S?q�@��?      �?              �?      �?(�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?      �?w&�1�L�?`ۛ:��?      �?                        6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @^Zq�$K�?ȖC�`��?      �?              �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?       @              @���@��?N#���?      �?              �?      �?$Zas �?              �?                                                              �?      �?      �?��N�Ա?ak�q�?      �?              �?        3~�ԓ��?      �?       @      �?               @       @               @       @              �?       @� Q�E��?�4ޫϹ�?      �?              �?        p�z2~��?      �?       @      �?       @               @       @       @       @      �?      �?      �?���>|�?2U�ui�?      �?              �?        ��RO�o�?      �?       @      �?                                       @                      �?       @J̖p���?,E�����?      �?      �?      �?      �?P�o�z2�?      �?       @      �?                       @       @       @       @      �?      �?      �?-?(�tN�?^a.�?      �?              �?        Zas �
�?      �?       @                       @       @               @       @      �?      �?       @A .��?�_�4�?                      �?      �?6���?              �?                               @       @       @       @       @      �?      �?�#�6���?T;���?�?              �?                ?���@��?      �?       @      �?                                               @              �?       @l	�Y �? zG�*�?      �?                        ���Vج?      �?              �?                                                              �?       @����e�?C��N.�?      �?                        $Zas �?      �?       @      �?                       @               @                      �?      �?j��|��?��	!��?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?�i)��X?      �?      �?                ���V؜?      �?       @      �?                       @               @                               @�5A .�?��<�?                      �?      �?6���?      �?       @      �?               @       @               @       @      �?      �?      �?s[ݧ���?�?���?              �?      �?      �?[as �
�?      �?              �?                       @       @       @       @              �?       @i�ae���?)#��\�?              �?      �?      �?ܥ���.�?              �?                       @                                      �?                �\d����?��<�?      �?                        ���V؜?      �?                       @                       @       @                      �?      �? .�c�?��V��?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                        ����'t�?;�0���?      �?                        v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?       @                ,1[�yj�?����?      �?              �?      �?      �?      �?       @      �?               @                       @              �?      �?       @+�oM��?�#�B�?      �?      �?                !�
���?      �?       @      �?                       @               @       @              �?       @�"X~PT�?W�A���?                              �?,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�d�Q�ϐ?�����?      �?                        �'�K=�?              �?                                       @                              �?       @P��*�?�S�Ȩ?      �?              �?              �?      �?       @      �?       @       @               @       @       @       @      �?      �?��-��?`{�D~�?      �?              �?        ��ۥ���?      �?       @                       @       @       @       @       @       @              �?T�@ʾ��?HPeB��?              �?                Zas �
�?      �?       @               @                                                      �?       @��7q��?�=/"Ӵ�?      �?              �?      �?p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @I`�:�?u�/����?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?              �?      @����[�? �<$3?                                �z2~���?      �?       @               @               @       @                              �?      @'���G��?#��^���?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?��sze��?              �?                              �?                       @               @                                      �?       @ͤ=����?`���|q?                                              �?                                                                                        ���"X~�?U�9��g?      �?                        �o�z2~�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                H���<�?���ƹ��?                      �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?���6�?>��Ϟ��?      �?                        F���@��?      �?       @      �?                               @       @       @              �?      @�$K!��?`[���?      �?              �?      �?�o�z2~�?      �?                       @       @       @       @       @       @       @               @J̖p���?=�B�80�?                      �?      �??���@��?      �?       @      �?               @                       @       @              �?       @�6��`�?�l�(��?                                �]�����?              �?                       @                       @       @              �?       @���7q�?R�����?      �?                        �@�6�?      �?              �?                                                              �?       @%�yO�0�?Y���?                                ��Vؼ?      �?       @      �?                                       @       @                       @�FR,?�?`@��ĸ?                      �?        6��9�?      �?       @      �?                       @                       @                      @h{����?^͜�ѻ�?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ��N�Ա?�e`���?                      �?        6��9�?      �?                                       @               @       @              �?      �?��9���?�kU�9��?      �?                        {2~�ԓ�?      �?                       @               @                       @                       @�����T�?��G��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?       @m+�oM�?�?Y�?      �?                        ���@��?              �?               @       @                                              �?      @SUUUUU�?����?                      �?        SO�o�z�?      �?       @                                                                      �?       @�����`�?���P�"�?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?       @t�ئ��?S�L�
�?                      �?        P�o�z2�?      �?       @      �?       @       @       @       @       @       @       @                P_W-��?^�q���?                      �?      �?�D+l$�?      �?       @      �?               @               @               @              �?        �Y;���?҅�)ǉ�?      �?                        {2~�ԓ�?      �?              �?               @               @               @      �?      �?      �?�=����?��b-��?      �?      �?                 �
���?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?E�(Ţe�?� L����?                      �?      �?      �?      �?              �?       @       @       @       @       @       @       @      �?        	�p���?���O�u�?                                ���V،?      �?              �?                                       @                      �?      @��<݌�?��'lߤ�?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @#w\I`ޓ?�Ր�,%?                                �@�6�?      �?       @      �?               @       @               @       @              �?       @7��+	�?�ަ�V�?      �?      �?      �?      �?$Zas �?      �?              �?       @               @       @               @      �?              �?J�hY7�?��PcK��?                      �?      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              @Y�)L�ْ?�����?      �?                      �?�o�z2~�?      �?                       @       @                                      �?                z����"�?��Y�̞�?      �?                      �?e�v�'��?      �?              �?       @       @               @       @       @      �?      �?       @[�KS}��?�C�K.r�?      �?      �?      �?        ��ۥ���?      �?       @      �?       @       @       @       @       @       @       @      �?        �c=kg��?��a$Y��?      �?                                      �?              �?                                                                      @D)-��?]v�{x?      �?              �?        >�]���?      �?       @      �?       @       @       @                              �?      �?       @�yjH��?���7�T�?                      �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        F��1��?{����?      �?                      �?�z2~���?      �?                       @                               @       @              �?      @�bѲ
n�?���\/�?      �?                                      �?       @      �?                       @               @       @              �?       @I�%��}�?@��F��?                      �?      �?F���@��?              �?               @                       @                                      @�'�F7��?�e`��?      �?              �?      �?�z2~���?      �?              �?       @                       @       @       @              �?       @䛌8j��?�k{S�?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?�p�t���?      �?              �?      �?Zas �
�?      �?                       @       @       @       @                       @      �?        F�Ɉ���?�����?      �?              �?      �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?����'t�?��_�?                      �?        P�o�z2�?      �?                               @               @       @               @                ٙ�ǰ2�?�����?                      �?        P�o�z2�?      �?       @      �?               @       @       @                       @              �?ʾ�����?�1�5k/�?                              �?���V،?      �?                       @                                       @              �?      �?q���Y�?m�_�R�?                                �'�K=�?      �?       @      �?                                                              �?      �?T�n�Wc�?�i��8�?                                �6��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?       @b��1��?E��t�?      �?      �?      �?        F���@��?      �?              �?                                                                        ��J��?�a_x��?                      �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?                      @1[�yj�?�w���?                      �?      �?��.�d��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @���C�?�w{�ɩ�?      �?                      �?              �?                       @                                                              @F�X�ڙ�?�V�φn?      �?              �?      �? �
���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�m��W�?t޶L\�?                      �?      �?p�z2~��?      �?                       @                       @                                       @�a/��?��c�7�?                                �ԓ�ۥ�?      �?       @               @               @       @       @       @      �?      �?      �?l�\d��?.�m�n��?      �?      �?                6��9�?      �?       @      �?       @                               @                      �?       @���l	�?�s�=�?                      �?        ,l$Za�?      �?       @      �?       @       @       @       @                              �?      �?{]�;x�?�H&X\��?      �?                        �D+l$�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @)g��1�?�S�o�?                                6��9�?              �?                               @                       @              �?      �?h�����?����?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�'�F7�?O���&?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?����T�?���5�?              �?                F���@��?      �?                               @                                              �?      @����?�/�B��?      �?              �?      �?(�K=�?      �?       @      �?       @       @                       @                      �?      �?�,���?�?�G�&���?                      �?        H���@��?      �?       @      �?       @                               @       @              �?      @#s�g�L�?�`��q��?      �?                        ���V،?      �?                       @       @                                              �?      @[ݧ����?'I���?      �?                        ?���@��?      �?                                                               @                       @����?�%�۔?      �?                        �z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?                       @)g��1�?٩w�!��?                      �?      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �j1v�?�(U9���?                                              �?              �?               @                                              �?       @�6��`��?5� ��kz?      �?                      �?�ԓ�ۥ�?      �?                                               @       @       @      �?      �?      @���q%�?;�E��I�?      �?                        ,l$Za�?      �?              �?               @               @       @       @                       @���?y4�?P�З�+�?      �?      �?      �?        �@�6�?      �?              �?                                                              �?       @��6���?��V/�?                                ���V،?      �?                               @                                              �?      �?��*��?����?      �?              �?        6��9�?      �?       @      �?                       @               @       @              �?       @P9��_��?@uc��?                      �?      �?�'�K=�?      �?              �?                       @               @       @              �?       @���.�?����h�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @����[�?>�G��U�?      �?              �?      �?�RO�o��?      �?                       @       @       @                               @                ����?"X�5%�?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      �?m+�oM�?|{��^�?      �?              �?        �K=��?      �?              �?       @       @                       @       @      �?      �?      �?�=�� Q�?�rC4��?      �?                      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @ś�8j��?��:��?      �?              �?      �?�o�z2~�?      �?               @      �?      �?      �?      �?      �?      �?       @                1[�yj�?�ۘx��?      �?      �?      �?      �?>�]���?      �?       @      �?       @               @               @       @      �?      �?        �o��z�?�7�^�S�?      �?              �?      �?6��9�?      �?                                       @               @                              @�
����?H|�$A�?      �?              �?      �?���@��?      �?       @      �?       @               @               @       @                      �?�<5���?���٧�?      �?                        F���@��?              �?               @               @                              �?              @�WH�%��?�Z�m�?      �?                        �]�����?      �?       @               @       @                                                       @^��C��?��r�3A�?      �?              �?        �K=��?      �?       @      �?               @                               @                      @5\.2�z�?���	��?      �?              �?        �'�K=�?      �?       @      �?               @       @                                      �?       @��H*��?)����?                      �?      �?��ۥ���?      �?       @      �?       @       @       @               @               @                ����e0�?d �S��?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?              �?        �'�F7�?���h��?                      �?        SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?                      �?E�(Ţe�?�k��a$�?      �?      �?      �?        Zas �
�?      �?       @      �?               @                                              �?       @:�X�?ҕ���
�?      �?              �?      �?      �?      �?       @      �?       @       @       @       @               @       @              �?e����I�?��V~���?                      �?      �?F���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        )g��1�?���Ъ��?      �?              �?        P�o�z2�?      �?       @      �?       @       @               @       @       @              �?       @����I{�?�Y���?      �?              �?        ��ۥ���?      �?       @      �?               @               @       @       @       @      �?      �?q���Y�?�x�� �?                      �?      �?6��9�?      �?              �?                                       @       @              �?       @5\.2�z�?�h2���?                      �?      �?��V��?      �?       @      �?       @               @       @       @       @       @               @�MF���?����p�?                      �?        �V�H�?      �?       @               @                                                               @}��j1�?������?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����'t�?\��Kd�w?      �?              �?        ?���@��?      �?       @      �?               @                       @       @              �?       @:'>���?RZ���?                      �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?�+Z��?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�U����|?�w�t2�?                      �?      �?	��V��?      �?                       @                       @                              �?      �?c9��?ޚL�
��?                                              �?                                       @                                      �?      @�%��f��?�|�:�m?                                �V�H�?      �?       @               @               @               @       @       @              @��.h�?3Ь�f�?                      �?      �?      �?      �?       @      �?       @       @                       @               @      �?        �	�p��?$�����?                      �?        $Zas �?      �?              �?       @               @       @       @       @      �?      �?      �?�oM���?��3�e�?      �?                                      �?                                                                                       @����e�?���W�g?                              �?�o�z2~�?      �?       @      �?                       @               @       @      �?      �?       @w\I`��?�\���?                                              �?                                                               @              �?       @��s��2�?�#h�q?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?޳J�6�?                      �?      �?�@�6�?      �?       @                                       @               @              �?       @q����?�Tt�T�?      �?                        �ԓ�ۥ�?              �?                       @       @                                      �?      �?�I�:Bl�?�%xH+�?      �?      �?                �]�����?      �?       @      �?                                       @       @              �?       @�N����?\%�|�?                                ���V؜?      �?       @                                       @       @                               @q��3��?�Ř�\�?      �?              �?      �?F���@��?              �?               @                       @                              �?       @ئ�N��?UҶ��ƞ?      �?      �?      �?      �?v�'�K�?      �?       @               @       @       @       @       @               @              �?)�tN|x�?BK����?      �?      �?                p�z2~��?      �?              �?       @                                       @                      @%K!�i�?n۶m۶�?                                      �?      �?              �?       @       @       @       @       @       @       @      �?       @Ͽk�.�?*k?i�?                      �?      �?      �?      �?              �?       @       @       @       @       @       @       @      �?      �?�x��?�`�~��?                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @                �%��}�?�H݇V�?                                Zas �
�?      �?       @      �?       @       @       @       @       @       @      �?      �?      @Z.2�z��?�2[�Y��?      �?              �?        ��RO�o�?      �?       @                                       @       @                      �?      �?�S�@��?+Iov9a�?      �?                      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?��q�S~�?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?                       @����'t�?�G�O��?                      �?      �??���@��?      �?       @                                                                              @���f���?c0|���?      �?      �?      �?        F���@��?      �?       @      �?                                                              �?       @̖p���?@*-���?      �?                        �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @                O�)���?Ge�g�?      �?                                      �?                                                                              �?      @�=�� �?t�Y=�h?                                �z2~���?      �?                               @               @                              �?       @����?��voǲ?                      �?      �?	��V��?      �?       @      �?       @               @               @       @              �?       @3��x�]�?	��uy�?                                F���@��?      �?                                       @       @               @                        8j��^�?N8�?a��?                      �?      �?���Vج?              �?                       @                                              �?       @�e0
84�? s���?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @1[�yj�?؄�3��(?      �?                        �z2~���?      �?       @      �?                       @       @       @       @              �?      @�#�d�Q�?���q�?                      �?      �?$Zas �?      �?       @       @      �?      �?      �?      �?      �?      �?              �?        <݌S��?�yr(ެ?                      �?      �?      �?      �?       @      �?       @       @               @                       @      �?        ����?���*�?                                ?���@��?      �?       @      �?                                                                       @k� 6\.�?�>�]ݢ?              �?      �?        ��RO�o�?      �?              �?       @                                                      �?        """"""�?X�F�28�?      �?      �?                �'�K=�?      �?              �?       @                       @       @       @                      �?��'t �?���i�?      �?              �?        (�K=�?      �?       @      �?       @       @               @                       @      �?      �?A��~5�?iX�=	�?              �?                F���@��?      �?                               @       @               @                      �?       @Ň7�B��?�(m�	�?      �?                        �D+l$�?      �?       @      �?               @       @       @       @       @              �?       @1�z�Τ�?���^�?      �?              �?      �?��RO�o�?      �?       @               @                       @               @                       @�?~�tт!�?                      �?      �?Zas �
�?      �?              �?       @               @               @       @                        ��S�@�?�`Q�6�?                                ���V،?      �?       @      �?                                                              �?       @x�ӥ�>�?��Z�m�?      �?              �?        ��RO�o�?      �?                                               @                                        d��ht�?�)�M�?                                ��ۥ���?      �?       @                               @                              �?               @ͤ=����?}1��#f�?                      �?      �?v�'�K�?      �?       @               @       @       @       @       @       @       @              �?8�B�]��?�!d&��?                                �K=��?              �?                               @       @       @       @              �?      �?��q
Sb�?��b�8K�?      �?              �?      �?      �?      �?       @               @                                               @                ��W��?F�F��G�?      �?                        ���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �j1v�?C#X�h`�?                      �?      �?F���@��?      �?                       @               @                       @              �?      @�^!ї�?W5=Dђ�?                                ���V،?      �?                                                                              �?      @ui��|��?�iN�Y��?                      �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @                E�(Ţe�?�K��C�?      �?      �?      �?                      �?              �?                                                                      @�9�፿�?�h�l��x?      �?              �?        ���V؜?      �?              �?                                                              �?       @p�l�?��*�t�?              �?                6��9�?      �?       @      �?       @       @                       @       @              �?        ���-�?�p)-��?                      �?        ���@��?      �?       @      �?       @               @               @       @      �?      �?      @A���Kn�?��*�@�?      �?                      �?v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?8�]�FR�?#�ۦw�?                      �?        ��RO�o�?      �?       @      �?               @       @       @       @       @      �?      �?        �}��?Ð�4b�?      �?                        ���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?����[�?*�r��?                                �@�6�?      �?                                               @       @       @                      @}�?^��?FZ(	Y�?      �?      �?                ���.�d�?      �?       @      �?                       @       @       @       @      �?               @1@�bѲ�?M�G5���?                      �?        >�]���?      �?              �?                       @       @       @       @              �?       @]d�����?�,�[���?                      �?      �?e�v�'��?      �?       @      �?       @       @                       @       @              �?        �����U�?�]|9��?      �?                        �ԓ�ۥ�?              �?               @               @                                              @��<݌�?����g�?      �?                      �?                      �?                                                                               @��w����?�b≋F?      �?              �?      �?���@��?      �?              �?               @       @       @       @       @      �?      �?        �p���?ع�(7D�?      �?                        ���V؜?      �?                                                       @                              @�a/��?������?      �?              �?      �??���@��?      �?                                                                                       @q%�yO��?�\kB+ӑ?      �?                        ���V،?      �?                                                                                        ~PT���?��_ͅ?      �?                      �?�ԓ�ۥ�?      �?              �?                       @               @              �?      �?       @Ͽk�.M�?wc^L!>�?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?�J%,h�?      �?                      �??���@��?      �?                       @                                                      �?       @��r�9��?�+Z��?                      �?      �?��RO�o�?      �?              �?       @                                                              @�u�b���?��]���?                                �@�6�?      �?       @      �?                                                              �?       @��x��?:Z�F�2�?      �?              �?      �?�'�K=�?      �?                                                                      �?      �?      @I`�:�?��VJM�?      �?                        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @h��2�?I�Mk'��?                      �?      �?�@�6�?      �?                               @               @               @      �?      �?        ��C��?o�8�*�?                              �?Zas �
�?      �?       @      �?                               @                      �?      �?      �?�?^���?�b��e�?                                                      �?                                                                      �?      @�j1v�?��Ub�G?      �?                        �@�6�?      �?              �?               @                                              �?      @�8�)1[�?xag��	�?                      �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�'�F7�?	��lR�?      �?              �?      �?3~�ԓ��?      �?       @      �?               @                               @      �?      �?       @Q��'�F�?��	��7�?                              �?!�
���?              �?               @               @       @       @       @      �?                mu����?U$�ڕ�?                      �?      �?              �?                                                                              �?        ��J��?�3�
'h?                                              �?       @                                                                      �?       @9�WH�?(���m?      �?                        v�'�K�?      �?                       @       @                                      �?      �?      @R��'�F�?1K���t�?                      �?      �?��.�d��?      �?              �?               @       @       @                                        ��H*��?>��
M�?      �?              �?      �?��V��?      �?       @                       @       @       @       @       @       @      �?        T�@ʾ��?��'��?              �?      �?        ���V؜?      �?              �?                                       @                      �?       @g��}���?1y���@�?                      �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?t+�oM�?N�����?                                ��RO�o�?      �?                       @       @                                              �?      @?(�tN|�?��G#�?      �?                        ���V،?      �?                                                                              �?      �?*g���?+T�ʟ?                                SO�o�z�?      �?                       @       @       @       @               @      �?              �?Q�E�*��?>���3�?      �?              �?      �?p�z2~��?      �?                       @               @                              �?      �?      �?��s��2�?ΡBY�3�?                      �?        >�]���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�c=kgҮ? �繫[�?      �?              �?      �?���@��?      �?       @                               @                              �?                ]!ї�V�?�o�8�*�?      �?      �?      �?        �D+l$�?              �?                       @                       @       @              �?       @�����`�?b���t��?      �?              �?        �'�K=�?              �?                                               @       @              �?       @���G���?al� g�?      �?                         �
���?      �?              �?               @                                      �?                ���I�:�?po��Ǉ�?                      �?        ��ۥ���?      �?       @               @       @       @       @       @       @       @                ~��j1�? �sjo�?                                Zas �
�?      �?       @                                                       @              �?        �U�����?��m�P��?      �?                        P�o�z2�?      �?       @               @       @       @                       @      �?              �?ï�Dz��?�[��<A�?      �?              �?        p�z2~��?      �?              �?       @                       @               @              �?       @O��b��?�k-|/�?      �?      �?      �?      �?p�z2~��?      �?       @      �?       @                                                      �?       @��*��?�u��v)�?                                �K=��?      �?              �?               @                                              �?      �?U:'>��?��3��?      �?                        {2~�ԓ�?      �?                       @       @               @                              �?      @��+	��?>�i�?      �?              �?      �?(�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @���6�?b���9�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @                F��1��?�>n΂�?                                �]�����?              �?                               @               @       @              �?       @F�X�ڙ�?+㇔&�?              �?      �?        �z2~���?      �?                       @               @       @       @       @      �?      �?       @��.h�?r����S�?                      �?        p�z2~��?      �?              �?                       @                       @              �?       @ J�hY�?N�'�0��?                                ���V،?      �?                       @                               @       @              �?       @L�*g��?���E�?      �?              �?      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?              @8�]�FR�?|�9G��?      �?      �?                6��9�?      �?              �?               @                                              �?       @O�0@�b�?`Ԋ;�ɳ?                      �?      �?�@�6�?      �?                                                                                      @�RG�mZ�?k��z�?      �?                        �@�6�?      �?       @      �?                               @               @              �?        ~��j1�?�8���?      �?              �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?ò
n�ͭ?-s���W�?      �?              �?      �?,l$Za�?              �?                               @       @       @       @      �?      �?       @����?�v�.��?      �?      �?                H���@��?      �?       @      �?               @                       @                      �?       @�����?�'w7��?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @��N�ԑ?q�w@o�?                                              �?              �?                                                              �?       @cX�~k��?EF�=?x?              �?                              �?              �?                                                              �?       @f��	��?�C�"J�x?      �?                        �]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�'�F7�?y!.�x��?      �?              �?      �?{2~�ԓ�?              �?                       @       @       @       @       @      �?              @�5\.2��?-�˕���?      �?      �?      �?        �D+l$�?      �?              �?               @       @                                      �?      @��<݌�?9K�T�?      �?              �?        �'�K=�?      �?                       @       @               @                       @      �?       @<�RG�m�?��ЏUW�?              �?                �RO�o��?      �?       @      �?       @                               @       @      �?      �?        �)1[�y�?m;{c���?                      �?      �?�ԓ�ۥ�?      �?                                                       @                              @ae��	�?G�Zln�?      �?                      �?�@�6�?      �?                       @       @       @               @              �?              @��6���?����<�?      �?                                      �?                                                               @                      @.������?���$�^q?      �?                        ��RO�o�?      �?       @                                                                              @}5&���?������?      �?              �?      �?v�'�K�?              �?                               @       @       @       @       @                �5A .�?79V$��?      �?      �?                �'�K=�?      �?       @      �?       @                       @               @       @               @���e0
�?X&s���?                      �?        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�X����?��nh:q?                                ���.�d�?      �?       @      �?                       @               @       @      �?      �?      �?��_���?G��hX�?      �?      �?                �D+l$�?      �?                       @       @                       @       @              �?       @F��s��?���0��?                                $Zas �?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?,1[�yj�?�����?                                Zas �
�?      �?                       @                                                      �?       @��"X~P�?hGEyI��?      �?                                              �?                                       @                                      @=Q�s�û?�	�+Z�S?      �?              �?      �?��V��?      �?       @               @       @                               @       @      �?      @���U�?ת�sze�?                                6��9�?      �?       @      �?                                                              �?      @�ئ�N�?����h�?                      �?      �?�@�6�?              �?               @               @               @       @      �?      �?       @ae��	�?<Q~���?      �?                                      �?              �?                                                                       @��j1v�?��7J-x?                      �?        �z2~���?      �?                                               @       @              �?                ٴ��I��?Ҷ��ƞ�?                      �?      �?�o�z2~�?      �?                       @               @                              �?              �?�`ph>�?���yr(�?                      �?      �?�K=��?      �?       @      �?               @       @       @       @       @      �?      �?      �?o��R��?޳J�6�?                                ��V��?      �?       @               @                       @                      �?               @���?y4�?�(u%ސ�?      �?              �?              �?      �?       @      �?               @       @       @       @       @       @      �?       @;�X��?����o�?      �?      �?      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        �S�@��?���SP2�?                      �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @��N�ԑ?em���?      �?              �?              �?      �?       @               @       @       @       @       @       @       @      �?      �?���@���?�%��Js�?      �?              �?        (�K=�?      �?              �?       @       @       @       @       @       @      �?      �?        �x��?��Z���?                      �?      �?��V��?      �?                       @       @       @                              �?      �?      @�������?:�첚�?      �?      �?      �?        �'�K=�?      �?       @      �?               @       @                       @              �?        Ž�,u��?��p��?      �?              �?        >�]���?      �?       @      �?       @                               @       @      �?      �?       @���?y4�?N
���K�?                                F���@��?      �?              �?               @       @                                      �?       @�b��!�?���Æ��?      �?      �?                �'�K=�?      �?       @      �?                                                                       @�B�]�F�?�fc���?                                F���@��?      �?              �?               @       @                                      �?       @�I�:Bl�?���L$�?                                              �?              �?                                                                       @J`�:�?�ͺ�ʏw?      �?                        �]�����?      �?       @      �?       @                               @       @              �?        �^<��u�?�v�.��?                                {2~�ԓ�?      �?              �?               @                                                      �?	�{B��?]�]����?      �?      �?      �?        �V�H�?              �?                       @       @       @       @       @      �?      �?        Ήo���?��`|���?      �?              �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @b��1��?��̈́y�?      �?                        ��Vؼ?      �?              �?                               @       @       @              �?        �	�p��?2;Mx[�?              �?      �?        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        n��W�?�탃�`�?      �?              �?      �?�ԓ�ۥ�?      �?              �?                               @               @              �?       @����q�?L;E��`�?      �?              �?      �?      �?      �?              �?       @       @               @       @       @       @                �����?���s	�?                      �?      �?�'�K=�?      �?                               @       @       @       @       @                        ��x��?|���{��?      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�፿Po�?fQ0���?      �?              �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�፿Po�?\�TQ��?                      �?              �?      �?       @      �?               @       @       @       @       @      �?      �?        ���\��?�DX�?|�?                                �D+l$�?      �?                       @       @                                              �?        ��W��?`�qpT�?      �?                        H���@��?      �?       @      �?               @               @       @       @      �?      �?        �S��%�?gQ���?                      �?        ���V،?      �?              �?       @                       @                              �?       @��̱���?�BcĔ?                                ���V؜?      �?       @      �?                                                              �?      �?��8j��?:)��Ý?      �?              �?      �?H���@��?      �?       @      �?                       @               @       @              �?       @!ї�V��?=1,��?                                ��RO�o�?      �?              �?                                                              �?      �?������?����q�?                                �6��?      �?       @      �?                       @       @       @       @              �?       @��8�)1�?~ z$Q�?      �?                              �?      �?       @               @       @       @       @       @       @       @                ��ds��?�sg����?              �?      �?              �?      �?       @      �?       @       @                       @       @      �?      �?        �~k� 6�?5�b��G�?      �?                                      �?       @      �?                                                              �?       @��8j��?g1'+<�z?      �?              �?      �?���.�d�?      �?       @      �?               @       @       @       @       @       @      �?      �?m�\d���?}u�/���?      �?              �?      �?6��9�?      �?                               @                                      �?              @B�/����?2X����?                              �?�z2~���?      �?       @      �?                                                              �?       @yO�0@��?�IGӹ?                              �?�z2~���?      �?       @      �?               @       @               @       @              �?       @���_���?7͉2k��?                      �?      �?��.�d��?      �?              �?       @               @               @       @      �?               @��'t �?k�h=�K�?              �?                >�]���?      �?       @      �?               @       @               @       @      �?      �?        �:Blӊ�?ψwG�?                      �?      �?�D+l$�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @n��W�?~|a�?                                $Zas �?      �?                               @                       @              �?      �?      �?,ZV���?��z�J�?      �?                                      �?                                                                              �?        ����7�?tO���h?      �?      �?                ���V،?      �?              �?               @                                              �?       @�6��`��?�*Œ�R�?                                ���V،?      �?       @                                       @                              �?      @��ǰ2��?��|8�?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                        �X����?����?      �?              �?        v�'�K�?      �?       @      �?               @       @                       @      �?               @�������?����~�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?E�(Ţe�?��ߧ��?      �?              �?        �'�K=�?      �?       @      �?       @       @       @       @       @                      �?       @�L�5A �?��|D���?      �?              �?      �?3~�ԓ��?      �?       @      �?       @                               @       @              �?      �?Q�����?5��0��?      �?              �?      �?v�'�K�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @F��1��?���\���?              �?      �?        ���V؜?      �?              �?                               @       @                      �?      @��J��?��Y
`�?      �?                        �@�6�?      �?              �?               @               @       @       @       @      �?      �?�p����?r��z�?      �?              �?        [as �
�?      �?                                       @       @               @              �?      �?�w�ӥ��?���5��?      �?      �?      �?        P�o�z2�?      �?       @      �?                       @                                      �?      �?���!���?���$Б�?              �?                              �?              �?                                       @                      �?       @��.h�?����T�|?      �?              �?        ��Vؼ?      �?                       @       @               @       @                      �?      @� �;�$�?���.���?                      �?      �?P�o�z2�?      �?       @               @       @       @       @               @      �?      �?       @��I{+�?���ܟ�?              �?      �?        ��ۥ���?      �?              �?               @       @               @       @       @      �?       @�O�n��?4��Ki��?      �?              �?      �?�K=��?      �?              �?                       @               @                      �?      @
Sb����?�UAZ�?                                p�z2~��?      �?                       @                       @                                      �?�Gm?C�?����?                                ܥ���.�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �??�]�FR�?,�x���?                                F���@��?      �?       @      �?                                                                      @���6�?��W�J�?                      �?        �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?                       @�bѲ
n�?�/�W~�?                              �?              �?                                                                                      @��}�ɣ�?��f�<�i?                      �?        ���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @<݌S��?x<��?      �?      �?                ���@��?      �?       @      �?                                       @       @              �?       @��.h#��?xX!�x��?      �?      �?      �?        ��ۥ���?      �?       @      �?       @       @       @       @                      �?      �?       @:Blӊ{�?�EF�=?�?                      �?        ��V��?      �?       @      �?       @               @               @       @              �?       @)���G��?Dtb�v�?                                $Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @              @^��Z��?w��?      �?              �?        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        8�]�FR�?G����?      �?              �?        �D+l$�?      �?                                       @                                      �?      @��e0
8�?���[Ӂ�?                                6��9�?              �?                                       @                                      �?*��:]�?e�[_:4�?                      �?      �?�'�K=�?      �?       @      �?               @                       @       @              �?       @S}䛌8�?�n����?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�፿Po�?@}m[&?      �?              �?      �?              �?       @      �?                                                              �?       @v���?�{�Sz?              �?                ���V،?      �?       @      �?               @                               @                       @���¯�?�b�B�ܐ?      �?                        >�]���?      �?       @      �?       @       @                                              �?       @݌S���?���c�?      �?              �?                      �?              �?                               @       @                      �?       @y4��0�?/̀�1?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?              �?       @nC��x�?M�Haw�?      �?                      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?                      �?�U�����?b�/��?      �?      �?      �?        p�z2~��?              �?               @                                       @                        R�&#��?���i6#�?      �?                        	��V��?      �?              �?                       @                                      �?       @=݌S��?d�+��?      �?                        ���Vج?      �?              �?                       @               @       @                        ӊ{'Y��?�f��?                                              �?               @      �?      �?      �?      �?      �?      �?                      �?8�]�FR�?����d!?      �?                        !�
���?      �?       @               @       @       @       @       @              �?      �?      �?�b��!�?��,�zU�?      �?                      �?�@�6�?      �?       @       @      �?      �?      �?      �?      �?      �?                      @�bѲ
n�?��:}�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                        #w\I`ޓ?�Ր�,%?      �?                                      �?       @      �?                                       @                      �?      @0��m$�?���%�?                              �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�፿Po�?���2�>r?      �?                        �z2~���?      �?       @      �?                       @               @                      �?       @�r�9ֳ�?�E�����?                      �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        #w\I`ޓ?�|�#��?                      �?      �?(�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @���Z��?m�w{���?              �?      �?              �?      �?       @      �?               @       @               @       @      �?      �?      �?�b�V��?D���?                      �?      �?$Zas �?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?��O��?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?t+�oM�?G&X\��?      �?                      �?���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @]����`�?6�4$�k?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ��Po��?���D�?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                      @���C�?/�F��G�?                                p�z2~��?      �?       @               @       @               @               @       @              @��#�d��?3H���?      �?                        [as �
�?      �?       @      �?               @       @               @       @      �?      �?       @Ţe� �?WDh���?                                �'�K=�?      �?              �?               @                       @                      �?        � �;��?��W�i�?      �?                                      �?                       @                                                               @{������?ҏ�;�k?      �?              �?      �?v�'�K�?      �?                       @       @       @       @       @              �?      �?       @��8j��?����q�?      �?                        �z2~���?      �?       @                               @               @       @                        F��s��?���U�?                                e�v�'��?      �?       @      �?               @                       @       @       @      �?        ��.h#�?�[Z���?                      �?      �?$Zas �?      �?       @      �?               @       @       @                      �?      �?       @�r�9ֳ�?�qM�F��?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @�'�F7�?wՐ�,e?                              �? �
���?              �?                               @                                      �?      @��Ͽk�?����?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?      �??�bѲ
�?���`��?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�U�����?��)~kw?      �?      �?      �?      �?6���?      �?       @      �?       @       @               @                      �?      �?        t3NaJ��?0�#���?      �?                      �?              �?              �?                                       @       @              �?       @�
n���?	���?      �?                      �?�z2~���?              �?               @       @               @                      �?                �U�����?�P�txn�?      �?                      �?              �?                       @       @               @               @              �?        ��J��?d�g$�ix?                      �?        P�o�z2�?      �?       @      �?                       @               @               @      �?        ��7q��? 7gA���?                                3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?                        �d�Q�ϐ?z9�=7�?                                ?���@��?      �?                                                                                      @Z��r�?O�mG�Z�?                              �?�]�����?      �?                       @       @                               @              �?       @H���<�?z7	t$�?      �?              �?        �ԓ�ۥ�?      �?       @      �?                                                              �?       @""""""�?Hz��	��?      �?              �?              �?      �?       @      �?       @               @       @       @       @       @      �?      �?V�ߚ ��?�e�U\�?      �?              �?      �?                      �?                       @                                                       @FaJ̖p�?�"!��U?      �?      �?      �?      �?p�z2~��?      �?              �?               @                       @              �?      �?        Ô�-�<�?�i^���?      �?              �?      �?���@��?      �?                       @                       @       @       @      �?               @���I�:�?K¥�H��?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?              �?      �?����[�?/(;p&k$?      �?                        �D+l$�?      �?       @               @                                       @              �?      @F��s�?�������?      �?                        ���Vج?              �?               @               @       @                                      @2&����?�y|�.�?                      �?        SO�o�z�?      �?       @               @               @       @       @       @       @              �?����?s��<�?              �?                �ԓ�ۥ�?      �?       @      �?       @       @       @               @       @      �?      �?       @wAIE��?X��I$a�?                      �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?                      @,1[�yj�?MD�i3a�?                                p�z2~��?              �?               @       @               @                      �?              �?���vA�?�э^�I�?                                F���@��?      �?                       @       @       @                                               @�o��z�?+����Ѩ?                      �?      �?6��9�?      �?       @      �?                                               @                       @l�\d��?�}xK�θ?                                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?��۩9�?                                �D+l$�?      �?       @      �?               @       @       @       @       @      �?              �?{�D_r[�?3�ߺ�n�?      �?              �?        �'�K=�?      �?                       @                       @                                       @�yjH��?�K¥�H�?                      �?        ?���@��?      �?                       @       @                                                      @E�*�A6�?0�����?      �?              �?        ���@��?      �?               @      �?      �?      �?      �?      �?      �?       @               @-h#���?��Y
`�?                      �?                      �?                       @       @                                              �?      @5\.2�z�?oj��lp?      �?              �?        ��RO�o�?      �?              �?               @                       @       @      �?      �?        ��s��2�?d�����?      �?                        �z2~���?      �?                                               @       @              �?      �?       @�^<��u�?o.����?                      �?        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�d�Q�ϐ?�Y@z�yi?                              �?�'�K=�?              �?               @                                       @              �?       @����?M3�z�n�?      �?              �?        {2~�ԓ�?      �?       @      �?               @       @               @       @      �?      �?        �*g���?���2���?                                F���@��?              �?               @                                                      �?        I`�:�?�B�[,�?      �?              �?        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�፿Po�?�D[T���?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @���C�?	�O��B�?                                              �?              �?                                                              �?       @��w����?˲T dQx?                      �?      �?�V�H�?      �?              �?                       @       @               @      �?                9�WH�%�? �R�3&�?              �?                                      �?                                                                      �?      @���Y;�?�U
u�wJ?                      �?        Zas �
�?      �?       @      �?               @                       @       @              �?       @.�jL��?���!d�?      �?              �?        �@�6�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @\��r�?/�K���?      �?              �?        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�d�Q�ϐ?K�q�h��?                      �?      �?��.�d��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @����'t�?t���B�?                      �?      �?              �?       @      �?       @               @               @       @              �?       @��E�X��?��6��ă?      �?              �?        [as �
�?      �?                       @       @       @       @               @      �?      �?      �?���I�:�?6j#��?      �?                        �ԓ�ۥ�?      �?                                                       @                              @jL�*g�?���;k�?                                �K=��?      �?       @               @       @               @                      �?      �?      @ .�c�?���}��?      �?      �?      �?        ��RO�o�?      �?       @               @                       @                      �?      �?       @`J̖p��?��]�t��?      �?              �?      �?�K=��?      �?       @                               @               @       @      �?                ��a�(��?�c>`�2�?                                              �?              �?                       @                                               @�Y e��?�l��{3{?              �?                ���V،?      �?              �?                                                              �?       @3NaJ̖�?�=k�?      �?              �?      �?���@��?      �?       @      �?       @       @       @               @       @      �?      �?       @�1���?�A[����?              �?                ���@��?      �?       @      �?                       @       @       @       @              �?       @�e� ��?+D�6�?      �?                      �?��ۥ���?      �?              �?               @                       @       @              �?       @c9�W�?����6��?                                �@�6�?      �?       @      �?               @                       @                      �?       @�d�#��?6��|g��?                      �?        6���?      �?       @      �?       @       @               @       @       @       @      �?      �?�"s�g��?,U��*��?                                [as �
�?      �?       @      �?       @       @                       @       @                       @}䛌8j�?�d�}���?                                ���V،?      �?                                                                                       @O�0@�b�?޵�8�?      �?                        ���V،?      �?              �?       @                                                      �?       @����J�?w�"�?      �?              �?      �?6��9�?      �?       @      �?                               @       @       @      �?      �?       @��U�?|���l�?      �?                        ?���@��?      �?       @      �?               @                               @              �?       @�^!ї��?E�����?                                �@�6�?      �?                       @                       @                      �?      �?      @9�WH�%�?m6a�E��?      �?                                      �?                                                               @              �?      @�yjH��?6��pq?                      �?      �?��ۥ���?      �?       @      �?       @       @       @               @       @       @      �?        _���@��?@Fg\�8�?              �?      �?      �?p�z2~��?      �?              �?                       @               @       @       @      �?       @�Up�l��?OsA=���?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�%��}�?��N�%�?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?u��U�?                      �?      �?���V؜?              �?                       @                               @                      @~(Ţe�?'gض�j�?                                              �?                                                                                      @�7�B�]�?#��=�g?      �?              �?        ���Vج?      �?       @      �?               @                                              �?       @?^��C�?D���<�?                      �?        �
��V�?      �?       @      �?                       @                                      �?       @��s���?x�]t�d�?      �?                        ��V��?      �?       @      �?       @               @       @       @       @      �?      �?      �?�d�#�6�?E(�DkJ�?      �?              �?        �@�6�?      �?                                                       @                                9�WH�%�?e�}��W�?      �?                                      �?              �?                                                                       @�V�ߚ�?x c[�cx?      �?              �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?ś�8j��?ޚL�
��?      �?              �?      �?H���@��?      �?                               @       @                              �?              @B����?z�Y�(��?                      �?      �?�z2~���?              �?                       @                                                      @S�KS}�?�Lb�&�?      �?                        �ԓ�ۥ�?              �?                                                                              @qi��|��?ꑂ/�?      �?                      �?��RO�o�?      �?       @      �?                               @                              �?       @�?^���?��9
��?      �?                        6��9�?              �?                               @                                              @�1���?��uV��?      �?              �?        6��9�?      �?       @      �?                                       @                      �?       @����q�?oy��|�?      �?      �?                ,l$Za�?      �?              �?                       @                                               @��Po��?vZ���?      �?      �?                ���Vج?              �?                               @       @       @                              �?�'t J�?0�'Tn'�?                      �?      �?�
��V�?      �?       @      �?                               @               @      �?      �?       @��ǰ2��?
�Nvd�?                                F���@��?              �?                                                       @              �?       @l��4�u�?#vQ��>�?              �?      �?        H���@��?      �?       @               @                       @       @                      �?      �?>�/�Q�?ÍC���?      �?              �?      �?�@�6�?      �?       @               @                               @       @      �?      �?        �8�)1[�?߮�wٜ�?                      �?        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����`�?EK^T��?                      �?        �D+l$�?      �?       @      �?                       @       @       @                               @Τ=����?y���?      �?              �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?        �%��}�?Z��Ґ?      �?                        6��9�?      �?       @                                               @       @              �?      �?���8�)�?��H�?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                g�)L�ٲ?�`�Z��?                                �z2~���?      �?                               @                                              �?       @��r�9��?��{�b��?                      �?      �?�z2~���?      �?              �?       @       @               @                                      @a�:�?m7���T�?      �?      �?      �?      �?v�'�K�?      �?       @      �?       @       @       @       @       @       @      �?      �?       @�e0
84�?��_�p��?      �?      �?      �?        (�K=�?      �?       @      �?               @       @               @       @              �?       @%��}��?�=�M'�?      �?              �?      �?�D+l$�?      �?       @               @                                                      �?        �ߚ ��?�� 0�?                                ��ۥ���?      �?                       @       @       @       @               @      �?      �?      @x�ӥ�>�?ڳ����?      �?                        ���V،?      �?              �?                                       @                      �?       @�`�AQ��?���^d�?      �?              �?        ��V��?      �?       @               @       @       @               @                      �?        �RG�mZ�?3��c���?      �?              �?        �RO�o��?              �?                       @       @       @       @       @              �?        �
����?.���]Q�?      �?                                      �?       @      �?                                                              �?      @��N���?�o��b5z?      �?                      �?�D+l$�?      �?                               @       @               @              �?              �?F��s�?
z��w:�?      �?                        e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�U�����?�Ҟ>�?                      �?        F���@��?      �?                       @               @       @       @       @                        \�՘H�?�F�oʔ�?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?       @�����`�?�E͙(t?                      �?        �@�6�?      �?       @      �?                       @               @       @              �?       @�۴���?,�;諭?      �?                        �RO�o��?      �?       @      �?       @       @       @       @       @       @      �?      �?      �?8�፿P�?�*�,%��?      �?                         �
���?      �?              �?               @       @               @                               @�hY7��?�n�N��?      �?      �?      �?        �'�K=�?              �?                       @       @                       @              �?      @yjH���?]V.դ?                      �?      �?�ԓ�ۥ�?      �?                       @       @               @                      �?      �?      @�:Blӊ�?F;h����?                      �?        �V�H�?      �?                               @                       @       @              �?      �?%�yO�0�?��C�A�?                              �?�]�����?              �?                               @               @       @      �?      �?      �?5w\I`��?�H���?      �?                        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?n��W�?�APx�S�?      �?      �?                H���@��?      �?       @      �?               @       @               @       @                      @�<5���?�G~�}x�?                                6��9�?      �?                               @               @               @      �?              @@�MF��?�1��?��?      �?                        �'�K=�?      �?              �?                       @       @       @       @              �?      �?��w�ӥ�?i~vT���?                                6��9�?      �?                               @                                                       @��Kn���?w$��S�?      �?              �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @F��1��?*N߆*�?      �?              �?        �D+l$�?      �?       @      �?       @       @       @       @       @       @       @               @��`ph�?CF͙(�?              �?                �z2~���?      �?       @      �?                       @               @       @      �?      �?        w\I`��?�'1�f�?                                ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ]����`�?����Æ�?      �?      �?      �?        6���?      �?       @      �?               @                       @       @              �?       @i�ae���?o����F�?                      �?      �?F���@��?      �?                       @                       @                      �?                ^!ї��?j_Ugw'�?      �?                      �?v�'�K�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�k�.M��?}�θ�q�?      �?      �?      �?              �?      �?       @                               @               @       @       @      �?      �?ui��|��?=O%���?      �?                      �?                      �?                                                                      �?       @�bѲ
n�?��A%OF?                                H���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��w����?Ǒo^��?      �?              �?      �?	��V��?      �?       @                       @       @       @                              �?      @ �&#���?"�)v�B�?                      �?      �?(�K=�?              �?                       @       @       @       @       @      �?      �?        ��r��?&Ve��<�?      �?                        !�
���?      �?       @      �?                       @                                              �?M+�d��?_���1�?      �?              �?              �?      �?               @      �?      �?      �?      �?      �?      �?       @                �Y;���?�f�����?                                P�o�z2�?      �?       @               @                                                              @�ߚ ��?cv݊�?      �?              �?      �?�D+l$�?      �?       @      �?       @       @               @       @       @       @      �?      @aѲ
n��?m����"�?      �?                        �RO�o��?      �?                       @       @       @                               @               @�o��z�?ԝ����?      �?                      �?��Vؼ?      �?                                                       @                               @c9��?�X�|v�?                                ��Vؼ?      �?                       @       @                       @       @              �?       @�k�.M��?�f�[_:�?              �?                >�]���?      �?       @      �?               @       @               @       @                       @�:Blӊ�?�O����?                      �?        �]�����?      �?                               @       @                                      �?      @E�*�A6�?�V�"�?                                ܥ���.�?      �?       @                       @       @       @       @              �?      �?        ��Po��?q-��yO�?      �?                        ?���@��?      �?                                                                              �?      �?q%�yO��?g���M��?              �?      �?      �?��RO�o�?      �?       @      �?                                       @       @              �?       @'t J��?�(ƾ���?                                H���@��?              �?               @       @       @               @       @      �?               @���vA�?[��'�x�?                                �RO�o��?              �?               @               @                       @      �?      �?       @�r@��?���X�?                                3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?      �?                F��1��?�gl��?      �?                        p�z2~��?      �?       @      �?                                       @       @              �?       @=���&�?Ǹ���?                      �?      �?���V،?              �?                                                                      �?      @����T�?r�V�u�`?      �?                        ?���@��?      �?       @      �?       @                               @                               @�ߚ ��?��E�נ�?                                3~�ԓ��?      �?       @                       @                                              �?       @�
����?T���j�?      �?                        $Zas �?      �?       @      �?       @       @                       @       @              �?       @�]�FR�?�`ּ��?      �?              �?        (�K=�?      �?       @      �?       @       @       @               @               @      �?      �?E������?�C�j��?      �?      �?                e�v�'��?      �?       @      �?               @                               @              �?       @�^!ї��?,�S�F$�?                                 �
���?      �?                               @       @                                      �?      �?�`ph>�?O\����?      �?                        �o�z2~�?      �?       @      �?       @       @                               @      �?      �?        �)����??��0�?      �?                        �]�����?      �?       @      �?                                       @       @              �?      �?�<݌S�?�Hվ���?      �?                      �?���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @#w\I`ޓ?�0g�~?                      �?      �?�]�����?      �?                       @       @       @                                              @�#�d�Q�?������?              �?                �'�K=�?      �?       @      �?                                               @                       @��`�AQ�?����b��?      �?                        ��Vؼ?      �?                       @                       @               @                      @Ň7�B��?c5XwA�?                      �?      �?�K=��?      �?       @      �?       @               @       @       @       @       @      �?      �?���(���?ZX�S[�?                                                      �?                                                                                ��N�Ա?�c[�cH?                      �?        �D+l$�?      �?       @      �?       @       @       @       @               @      �?      �?      �?��I�:B�?��<���?                                3~�ԓ��?      �?       @      �?               @                       @       @       @                O����7�?p�$6�?                                e�v�'��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @���@��?c"�;
�?      �?                      �?3~�ԓ��?      �?       @                       @       @       @       @       @      �?              �?�ǰ2���?�J���N�?      �?                                      �?                               @                                                       @]<��u��?1��?n?                      �?      �?(�K=�?      �?       @               @                       @       @       @       @      �?        r�g�L��?��=��?                      �?      �?	��V��?      �?       @      �?                                               @              �?       @b�(Ţe�?��R,�)�?      �?                         �
���?      �?                       @                       @       @       @      �?                �N���?T������?      �?                        �o�z2~�?      �?       @      �?       @       @       @                                                j��|��?��Ys��?                      �?        �]�����?              �?               @                       @                                        Y�՘H�?:L����?      �?                        F���@��?      �?       @      �?                                               @              �?       @���w���?�=��-ű?                                �'�K=�?      �?       @      �?               @                       @       @              �?       @w\I`��?ק�T��?                                ���V،?      �?              �?       @               @                                      �?       @*L����?	R9���?                                              �?                                                                                      @�����9�?���W�i?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?              �??�TS��?                      �?      �?6���?      �?              �?       @       @                       @       @      �?              �?����?0K@��?                                �'�K=�?      �?       @                                               @       @      �?      �?      �?������?�_7r�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      �?nC��x�?��q�S~-?              �?                6��9�?      �?       @      �?                                       @       @              �?       @�Up�l��?<���eM�?                      �?      �?�o�z2~�?              �?               @       @               @       @               @                Y���d�?�?93q�?              �?      �?        ��ۥ���?      �?              �?       @       @       @       @       @       @       @      �?        
���O�?,v��$�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?_�<$3h?      �?                        �'�K=�?      �?       @                                               @                      �?       @��2�?>,*��?                                �ԓ�ۥ�?      �?       @      �?               @                       @                      �?      �?��,u���?�ZNy&H�?                                ���Vج?      �?              �?               @               @               @              �?       @�G�Ɉ��?�r�*�?                                              �?                                                                              �?       @��j1v�?�����g?      �?                        �z2~���?      �?                                                                              �?        �'t J�?ֽ�����?                                �D+l$�?      �?                       @       @       @       @       @              �?              �?�k�.M��?AN����?                                �z2~���?      �?       @      �?       @       @                               @      �?                ��C���?�W���U�?                      �?        ���V،?      �?              �?       @       @                       @                               @����?����I�?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?�x
JƓ?                                �
��V�?      �?                               @               @                                        �5A .�?;����"�?                                �K=��?      �?       @                                       @       @                              @I!�i��?�pL���?      �?                        F���@��?      �?       @       @      �?      �?      �?      �?      �?      �?                      @s�rv��?��{i�8�?      �?              �?      �?�z2~���?      �?                       @                       @                       @                �5A .�?��I���?                      �?        ��RO�o�?      �?       @               @       @       @                       @      �?                ]�;x��?'����,�?                                p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?qi��|��?������?                      �?        �
��V�?      �?       @      �?                       @       @       @       @              �?       @Y7���?���W[�?      �?              �?      �?�K=��?      �?                       @               @       @               @       @              @-h#���?I9��?      �?                        6��9�?      �?       @      �?               @                                                       @��*��?Ǯ�����?      �?                        p�z2~��?              �?               @                               @       @      �?      �?      @F�X�ڙ�?]-a����?                      �?      �?(�K=�?      �?       @      �?               @       @               @       @      �?      �?       @C��x�?�J@_�>�?      �?                        �'�K=�?      �?       @                                                                      �?       @}5&���?!�����?      �?              �?              �?      �?       @      �?               @       @               @       @       @      �?        Wc"=P9�?����?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @F��1��?�?��Ӎ?      �?              �?        ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @n��W�?�bk��?      �?              �?        (�K=�?      �?       @      �?       @       @       @       @       @       @      �?              �?�䶺O�?;��5[�?                                3~�ԓ��?      �?       @               @                               @       @      �?              @F��s��?��6&���?                                �'�K=�?      �?                       @               @       @                      �?              �?�Wc"=P�?����mW�?                                              �?              �?                                                              �?       @�c9�?o��W�w?      �?              �?      �?p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @n��W�?eCW�ڍ�?                      �?        ��ۥ���?      �?                               @       @       @       @       @       @      �?      �?�AQ�s��?��z`;��?      �?              �?      �?�@�6�?      �?       @               @       @       @               @                      �?      �?9ֳv&��?�!�0�?                      �?      �?(�K=�?      �?       @      �?               @       @       @       @       @       @      �?       @��|�G�?�P�KlS�?                      �?        F���@��?      �?       @      �?                                       @                      �?       @c"=P9��?j����?                      �?      �?Zas �
�?      �?       @      �?               @                       @       @              �?       @9�)1[��?SH���?      �?                        F���@��?      �?       @      �?               @                       @       @              �?       @!ї�V��?y@�;U�?      �?                                      �?              �?                                       @       @              �?       @O��b��?v�1/��?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @,1[�yj�?�3��o��?      �?                      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?� Co8X�?      �?              �?        	��V��?      �?       @      �?               @       @               @       @              �?       @a/���?���u�?                      �?      �?p�z2~��?              �?               @       @       @               @       @      �?               @��c�?��%���?      �?              �?      �?���V،?      �?       @               @                                                              @?(�tN|�?�LRd�?                                ?���@��?              �?               @               @                                              @SUUUUU�?hexSh��?      �?                        ?���@��?              �?               @       @               @                                      @�8j���?E���'�?      �?      �?      �?        ��V��?      �?       @      �?               @                       @       @              �?        S}䛌8�?���6�?                      �?      �?�RO�o��?              �?               @               @       @       @       @       @              �?G�%��}�?#g�`�?      �?                        �RO�o��?      �?       @      �?               @                       @                      �?        8�B�]��?�C��?                      �?      �?�z2~���?              �?                                       @                      �?              �?b��1��?����t��?                      �?        �@�6�?      �?       @      �?                                       @       @              �?       @��1��?6��P�?      �?      �?      �?        Zas �
�?      �?                       @       @                                              �?        �
n���?���ѷ?      �?                        �
��V�?      �?       @      �?               @                       @       @      �?               @:'>���?.-GB��?                      �?                      �?               @      �?      �?      �?      �?      �?      �?              �?      @����'t�?�>�!�+?                                �'�K=�?      �?              �?               @       @               @       @              �?       @;�RG�m�?<�+R?�?      �?                        H���@��?      �?       @      �?                                               @              �?       @y4��0�?��m����?      �?                        3~�ԓ��?      �?       @      �?                                               @              �?        o��4�u�?���ə��?              �?                ���V،?      �?       @      �?                                       @                      �?       @�}�m�?eb%��?      �?      �?                SO�o�z�?      �?       @      �?               @                                              �?        d��ht�?����Վ�?      �?              �?        p�z2~��?              �?                               @                                               @'���G��?�6��ĳ?                                �D+l$�?      �?       @      �?               @       @                                      �?       @ئ�N��?)ִ8�4�?      �?              �?      �?{2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?              �?        ���C�?"b/�v�?      �?              �?      �?(�K=�?              �?                       @       @       @       @       @      �?               @��E�X��?7�g�m�?              �?      �?                      �?       @      �?                       @               @       @              �?       @_���H�?��g��`�?              �?      �?        Zas �
�?      �?       @      �?       @       @       @       @                              �?      �?���.�?��ɼ7��?      �?      �?                ��ۥ���?      �?       @      �?               @               @       @       @       @      �?       @ճv&�1�?�D@w�?                                p�z2~��?      �?       @      �?       @                       @                              �?       @����?��PHY�?                                ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                        nC��x�?;�6���?      �?                        6��9�?      �?              �?               @       @                                      �?       @�rv��?�� ����?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @nC��x�?9��.��?      �?              �?        SO�o�z�?      �?       @               @                                              �?              �?�%��}�?�
E}�?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @#w\I`ޓ?�G�O���?      �?                        ��V��?              �?                       @                       @              �?      �?       @R�&#��?F����?      �?              �?      �?�
��V�?      �?              �?                       @               @                               @b�(Ţe�?�3�����?      �?              �?        	��V��?              �?               @               @                                              @�Po���?�Rj�t��?                                ,l$Za�?              �?                               @               @       @      �?      �?       @��*��?�ǟn���?                              �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?c�����?      �?      �?      �?        (�K=�?      �?       @               @       @       @       @       @       @       @      �?      �?��q
Sb�?1؈��7�?                                6��9�?      �?              �?       @                               @                      �?      @��a�(�?d�(�$�?              �?                �V�H�?      �?       @                               @       @               @      �?      �?      �?%�yO�0�?r)�B��?                                �D+l$�?      �?       @                       @       @               @              �?      �?      �?� �;�$�?�Z�����?                              �? �
���?              �?               @                       @               @                      @����U��?�_/���?                                �
��V�?      �?       @                                       @                              �?      �?]!ї�V�?1�+5��?                      �?      �?�D+l$�?      �?       @               @               @       @       @               @      �?      @0�	��?SR���?                                �'�K=�?      �?       @                                                                      �?      @d��ht�?{�ڇ��?      �?                        6��9�?      �?              �?                                                              �?      @3NaJ̖�?�u����?      �?      �?                ���.�d�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        n��W�?ɍ �j�?      �?              �?      �?�'�K=�?      �?                                                                                        �d�Q���?ITC���?      �?                      �??���@��?      �?       @      �?               @                       @       @              �?       @��6��?���;km�?      �?                                      �?                                                                                       @�����9�?���W�i?                                �'�K=�?      �?                       @       @               @                      �?                ��	�p�?��G����?      �?                      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @�%��}�?9��.��?                      �?        >�]���?      �?              �?       @               @                               @                ������?���S���?      �?                        ���V،?      �?              �?       @       @                       @       @                       @:'>���? a��;�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @E�(Ţe�? ��??      �?      �?                6��9�?      �?       @      �?                                       @       @              �?       @KS}䛌�?
s�����?                                �]�����?      �?              �?               @       @               @                      �?       @嶺O_�?|M"	�?              �?      �?        �o�z2~�?      �?                       @               @       @       @       @       @      �?      �?�`�AQ��?2���Z��?                      �?        �'�K=�?      �?              �?               @       @               @       @                       @�3i�ae�?	zb2X�?      �?      �?                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�'�F7�?�7$�_��?                              �?              �?              �?       @                                                      �?      @�Ɉ����?�ꖜ��y?                                ��ۥ���?      �?                       @       @       @       @       @              �?      �?      @�Y e��?'ʬA
�?      �?              �?      �?              �?              �?                                                              �?       @      �?�_���}w?                                �@�6�?      �?              �?                                                              �?      @o�Wc"=�?l�q䛧?      �?      �?      �?        �@�6�?      �?       @      �?       @               @                                      �?        x�����?���s	�?      �?              �?      �?[as �
�?              �?               @                       @                                        �������?�j<�WF�?                      �?        �@�6�?              �?               @                                                               @��2�?eX�=	�?      �?              �?      �?H���@��?              �?               @                                       @              �?       @ku����?�4Z��?      �?                      �?              �?       @      �?                       @               @       @              �?       @^��C��?}��m!�?      �?              �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @��N�ԑ?E-�<$�?      �?              �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        !�iŽ�?́��B�?      �?                        �@�6�?      �?              �?       @               @                                      �?        �?^���?s�A��?              �?                ?���@��?      �?       @      �?                                                              �?       @�@ʾ���?X)�*I�?      �?                        ��Vؼ?      �?              �?                                                              �?       @}�?^��?JHy�f�?                      �?        p�z2~��?      �?                       @               @               @              �?      �?      �?MaJ̖p�?����,�?              �?                ���Vج?      �?                       @       @               @                                      �?Ήo���?P��T�ʟ?                                �@�6�?      �?              �?       @       @       @       @               @              �?        ��	�p�?&;2E 5�?                      �?      �?6��9�?      �?       @      �?               @       @                       @              �?       @?(�tN|�?d6�����?                      �?      �?P�o�z2�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ,1[�yj�?R�\
���?      �?      �?      �?      �?���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ����T�?q`^����?      �?                                      �?              �?                                                              �?       @�l	�Y�?�-˽x?      �?              �?      �?>�]���?              �?               @       @               @       @              �?      �?      @�@��~�?k�+�*�?              �?      �?        p�z2~��?      �?       @               @       @       @                                      �?      �?�����T�?� [���?                                      �?      �?       @      �?               @       @       @       @       @       @      �?        �B�/��?>�ts���?              �?                �ԓ�ۥ�?      �?              �?                       @                       @              �?       @Ô�-�<�?[ł���?                      �?         �
���?      �?       @      �?               @                                                        ���Up�?�����?                                �'�K=�?              �?               @       @       @       @                      �?              @���G���?[�����?                      �?      �?Zas �
�?      �?       @      �?               @                                              �?      �?�`�AQ��?>�"�Ms�?                                �z2~���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @^��Z��?�=�t��?                      �?              �?      �?       @      �?               @       @       @       @       @      �?              �?��g{��?O�ñ�?                                              �?                                                                              �?       @�����9�?���W�i?      �?                              �?      �?       @      �?       @       @       @       @       @       @       @                s@���K�?T�<���?                      �?        �V�H�?              �?                                               @       @              �?       @�7�B�]�?L��	a�?      �?                                      �?                               @                                              �?       @ئ�N��?X2��3n?              �?                              �?       @      �?                                                              �?       @���q%�?��=1y?      �?              �?        P�o�z2�?      �?              �?               @               @       @       @      �?      �?       @��'t �?�`#�#��?      �?              �?        v�'�K�?      �?       @      �?               @               @       @       @      �?      �?       @�#�d�Q�?�Oˊ^_�?      �?                      �?�6��?      �?       @      �?               @                                              �?      @�yO�0@�?�[}/-�?      �?      �?      �?              �?      �?       @               @       @       @               @       @       @      �?      �?�W���?	�B��?      �?                        ��V��?      �?       @      �?       @                                              �?                ���U���?�4F�?      �?      �?                6��9�?      �?       @      �?               @                       @                      �?       @M���E�?(#�Ǘ��?              �?                �'�K=�?      �?              �?                                       @       @              �?       @�V�;�R�?�x(?�g�?      �?                        $Zas �?              �?                               @       @                      �?              @�.h#��?�~^��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @����[�?/(;p&k$?      �?              �?      �?6��9�?      �?                       @               @       @                      �?      �?      @����?X�*�!�?                      �?        (�K=�?              �?               @       @       @       @       @       @       @                ���>|�?��ع��?      �?              �?      �?���.�d�?      �?       @      �?                       @                       @      �?              �?���@���?�څ�{��?      �?      �?                              �?              �?                                                              �?       @����e�?M�$&�x?      �?                        3~�ԓ��?      �?       @      �?               @               @       @       @                       @��Ͽ�?�t�Y=��?                                �z2~���?      �?       @      �?                                       @       @              �?       @���.�?��?��X�?                      �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?                        �፿Po�?�yW��/�?              �?                H���@��?      �?       @      �?                       @                       @              �?      �?�
n���?.F����?              �?      �?        ���V؜?              �?                       @                                              �?       @_ph>׿?���E~?                      �?        �'�K=�?      �?       @      �?       @                               @       @              �?       @�p����?�^ۛ:�?                      �?      �?���V؜?              �?               @                                                              �?P��*�?��nh:�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @�U����|?�;�N���?                      �?              �?      �?       @               @       @       @       @       @       @       @      �?       @T��%��?}<a�&��?              �?                �z2~���?      �?              �?       @       @               @                              �?        1v�z�?���[��?                                              �?       @      �?                                               @                      @��H*��?�^,5�?                                ���V،?              �?                       @                       @       @                       @�>�MF�??3�z�n�?                      �?      �?�z2~���?      �?                       @       @       @       @                      �?      �?      @f��1��?����`�?      �?              �?        P�o�z2�?      �?       @               @       @       @       @       @       @       @      �?      �?�?y4��?�U4�?      �?              �?        �6��?      �?              �?       @       @                                              �?       @�ti��|�?N�-��?      �?      �?      �?        �ԓ�ۥ�?              �?                               @                              �?      �?      �?��Ͽk�?���x(?�?                      �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?                       @,1[�yj�?�_M좤�?      �?      �?                              �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?�^/��"?      �?                        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @���@��?��w��V�?                                �
��V�?      �?       @      �?       @               @                              �?      �?      �?~5&��?�����?                      �?        �'�K=�?      �?       @      �?               @       @       @       @       @      �?      �?        x�/���?�j�i��?                                F���@��?      �?       @      �?                                               @              �?       @l�\d��?�tU����?              �?      �?        ��ۥ���?      �?              �?               @       @                       @       @              �?[ݧ����?��w~��?      �?              �?        �K=��?      �?       @               @       @       @       @                       @              �?��=���?�qhف3�?      �?              �?        �ԓ�ۥ�?      �?       @      �?               @               @       @               @      �?      @c9��?���h��?      �?                        ?���@��?      �?       @                                       @               @                      @�*��?6��x�Ι?      �?                                      �?                                       @       @       @       @              �?       @���I�:�?�Ms��z?                                6��9�?      �?                                       @       @                                       @���@���?�ȸ��?      �?                        ��V��?      �?                               @       @               @                      �?      �?�w�ӥ��?�Rb�q�?                      �?      �?>�]���?      �?              �?                                       @       @      �?                �&#��~�?�	W�~F�?      �?              �?      �?��V��?      �?                               @       @       @       @       @       @              �?Po��T�?��E��?      �?                        �z2~���?      �?                               @                                              �?        ��*��?` �e���?      �?              �?      �?�@�6�?      �?                                       @               @                      �?        .��:]�?	^��ڠ�?                      �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        m+�oM�?1C�Lޣ�?      �?      �?      �?      �?P�o�z2�?      �?               @      �?      �?      �?      �?      �?      �?      �?                nC��x�?#�'�Y�?                                �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�፿Po�?���ݰ��?      �?              �?      �?�z2~���?              �?                       @               @                                      @���[��?�
"_m�?      �?              �?      �?>�]���?      �?       @      �?       @       @       @       @       @       @       @              @��*��?�E��.�?      �?                        ���Vج?      �?                                       @       @                                       @z����"�?�n���?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                        F��1��?^mT�Et�?                                �'�K=�?      �?              �?       @                               @                               @�a�(Ţ�?�kѥ�{�?      �?              �?      �?(�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?qi��|��?%E�r�)�?      �?              �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @m+�oM�?����E�?      �?                      �?��RO�o�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?����[�?�a��-��?                      �?                      �?              �?                                       @                      �?        d��ht�?����z�|?      �?              �?      �?�6��?      �?                       @               @       @       @       @       @              �?�����?��g?ʤ�?              �?      �?        $Zas �?      �?              �?       @       @                       @       @      �?              @u�4�G��?�ۃ�"��?                                H���@��?      �?                       @       @       @       @       @              �?              @j�����?!���V@�?      �?      �?                Zas �
�?              �?                       @                       @                      �?      @<�RG�m�?��U�$��?                                �@�6�?      �?                                                                              �?      @�d�Q���?s��]ʪ?                                �z2~���?              �?               @               @       @               @       @              @h#���?i�K���?      �?                        �@�6�?      �?              �?               @                                                       @S,ZV��?�d�}���?                      �?                      �?              �?                                       @                               @)���G�?��F�[|?      �?      �?                ��RO�o�?      �?       @      �?                                                              �?       @S,ZV��?Ir�g,�?      �?              �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?#w\I`ޓ?u5�9���?      �?      �?      �?        �@�6�?      �?              �?                       @               @       @              �?       @d�#�6��?�8��d�?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?.�r@�?"�:1z�?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����`�?�'�'�?      �?              �?      �?�@�6�?      �?              �?                                                              �?       @ї�V�i�?��|W�6�?      �?      �?                ��V��?      �?       @      �?       @               @       @       @       @       @      �?       @��Z�KS�?��,
��?      �?      �?                              �?                                                                                       @����7�?tO���h?      �?                        {2~�ԓ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @_����,�?����@7�?                      �?      �?���V،?      �?              �?                                                              �?       @�=�� �?hexSh��?                              �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?�k�*���?                      �?      �?$Zas �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        m+�oM�?����0��?                              �?F���@��?              �?               @                                                              @��Ͽk�?��<��?      �?                                              �?                                                       @                       @3\.2�z�?��)*`?              �?                              �?              �?                                                              �?       @o�Wc"=�?\��Kd�w?                      �?      �?��.�d��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ?�]�FR�?� |�?      �?      �?      �?        6��9�?      �?              �?               @       @       @       @                      �?      @�-�jL��?�\���	�?      �?                        �z2~���?      �?       @      �?                                       @       @                       @�0%fK�?��W[�?                      �?        $Zas �?      �?              �?                                                              �?        ї�V�i�?�m�ZNy�?      �?              �?      �?H���@��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�6��w�?����?                      �?      �?��ۥ���?              �?               @       @               @       @       @       @                �3i�ae�?)�+u�N�?                              �?                      �?                                                                              @�bѲ
n�?��A%OF?                                              �?               @      �?      �?      �?      �?      �?      �?                       @F��1��?��ֺ�?      �?                        �D+l$�?      �?       @                               @                               @              �?^!ї��?��z���?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?                        8�]�FR�?����d!?      �?                        ���.�d�?      �?       @               @       @       @       @       @              �?               @\�՘H�?퐷�@}�?                                �]�����?      �?              �?               @                               @              �?      @�H*���?�%�ׅ!�?      �?              �?        �V�H�?      �?                       @       @       @       @                       @              @��a/�?�Blk]�?      �?      �?      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?n��W�?j��s�'�?      �?              �?      �?�
��V�?      �?       @                       @                               @                       @ .�c�?�VHV:W�?                                SO�o�z�?      �?                                       @       @               @       @              �?��C��?B�w"�C�?                                ��RO�o�?              �?               @       @       @       @       @              �?      �?       @�����?ڪe��?      �?      �?      �?        �'�K=�?      �?       @      �?                       @               @       @              �?       @P9��_��?#�Ҟ�?                      �?      �?�]�����?      �?                                                       @                               @z����"�?�����Q�?      �?      �?                	��V��?      �?              �?               @       @               @       @              �?       @��:]��?��"2M��?      �?      �?      �?        �'�K=�?      �?       @      �?                                       @       @              �?       @�Gm?C�?I��<wu�?      �?                      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?ò
n�ͭ?���F}֨?      �?      �?                F���@��?      �?       @      �?                                                                      @*g���?�X����?              �?      �?        p�z2~��?      �?       @      �?                       @               @       @                       @�;�$0��?�1��u�?      �?              �?      �??���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�d�Q�ϐ?�G���W{?                      �?        ���.�d�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����'t�?Z���[��?      �?                        ,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?       @              @n��W�?�<���i�?      �?      �?                �z2~���?      �?                       @               @                       @      �?              �?+?(�tN�?} z�?      �?                        �z2~���?              �?               @       @               @       @                      �?        �������?y�\�V�?      �?              �?        [as �
�?      �?       @      �?               @       @               @                               @����C�?ߴ�$)�?                                $Zas �?              �?                       @       @       @                                        H���<�?!�/n�O�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      �?,1[�yj�?p�/
b7�?                                �
��V�?              �?                               @                                      �?      @eZq�$K�?�N &pͶ?                      �?      �?�@�6�?      �?              �?               @                                              �?        ��#�d��?�y�(��?              �?      �?        �]�����?      �?       @               @       @               @                              �?      @-����?3��j�!�?                      �?      �?�ԓ�ۥ�?              �?               @                       @       @               @      �?      �?�@ʾ���?";��zE�?      �?              �?      �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              @^��Z��?g��,��?      �?                                      �?                                               @                                      �?}5&���?����T�l?      �?              �?      �?�]�����?      �?       @      �?       @               @       @                      �?      �?      �?�`ph>�?ad����?      �?                        H���@��?      �?       @                                       @       @               @      �?        [�<��?oy��|�?      �?                        ��RO�o�?      �?              �?                                                              �?      @b����,�?��8�5�?                                ��RO�o�?      �?              �?                                       @       @              �?      @�hY7��?ZNy&Hf�?                                F���@��?      �?              �?               @                       @       @      �?      �?      @z����"�?�>?(�?                                �RO�o��?      �?              �?               @       @               @       @       @      �?       @�p����?�:�R��?      �?              �?      �?���.�d�?              �?               @               @       @       @       @       @      �?        `J̖p��?���B�?      �?                                      �?              �?                                       @                      �?       @����[�?R�3.z|?      �?                        3~�ԓ��?      �?              �?                               @       @       @              �?       @Aʾ����?��_�?                      �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @                ���C�?�zj�,�?                                �6��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�'�F7�?|�Ѡe�?                                �ԓ�ۥ�?      �?                       @       @       @                                               @�!�����?�nE��?                      �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @              @�5A .�?|Ck�+�?                      �?      �?p�z2~��?              �?               @       @       @       @               @       @      �?      @1���?���/��?      �?              �?      �?�ԓ�ۥ�?      �?                                       @                       @                       @�Y;���?O�c���?      �?      �?      �?        ���V،?      �?       @      �?                                       @                      �?      @�������?n��
�@�?      �?              �?      �?SO�o�z�?      �?                       @       @                                                      @,u�ئ�?�����?      �?                        �6��?      �?       @      �?               @       @                       @              �?      �?{]�;x�?�1/��?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @                �d�Q�ϐ?Rke����?      �?                        ���V؜?      �?                                                                                      @B�]�FR�?��a�?                                              �?       @      �?               @                                              �?      @ZV����?n�CT}?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?�b/��?                                                      �?                                               @                      �?       @Sb����?V�φ^?      �?                        ��Vؼ?              �?               @       @       @                              �?              @¢e� �?�"R9�?      �?                        $Zas �?      �?       @      �?                               @       @       @              �?      @��r��?���&��?      �?      �?                �@�6�?      �?              �?                       @               @       @              �?        fK8O��?Nn��?              �?      �?        �]�����?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                Rp�l?Q;�m,P�?      �?              �?      �?H���@��?      �?                       @                       @                                       @����?�_�3d��?                      �?        F���@��?      �?                       @                                                      �?         e��h�?w\�.}ޣ?                      �?        $Zas �?              �?               @               @               @       @                       @������?�$�hh��?      �?              �?        ���Vج?              �?                                                                      �?       @�?UT��H�?              �?      �?        ��V��?      �?       @      �?               @       @               @       @      �?      �?       @s��2�?j�V�A��?      �?                        $Zas �?      �?              �?       @       @       @       @       @       @              �?        -�<5��?0�ۃ�"�?      �?              �?      �?	��V��?      �?              �?                                       @                               @B�/����?�B��i�?      �?              �?        	��V��?      �?                       @       @                               @      �?              @1�z�Τ�?	���?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?      �?              @���C�?ݘ<$3(?      �?                        $Zas �?      �?                               @                                              �?      @��>|]�?��i>���?                      �?        6��9�?              �?               @                       @       @               @               @�'t J�?�����@�?      �?              �?        Zas �
�?      �?       @                       @       @               @       @       @                m$���?�\P�$�?      �?                      �?$Zas �?              �?                               @       @       @       @      �?                ؋�ߵN�?R�	��?                                �K=��?      �?                       @       @               @                      �?              �?����?��q�?              �?      �?        �ԓ�ۥ�?      �?       @      �?                       @               @       @                        mu����?㇔&�[�?                                ���.�d�?      �?       @               @       @       @       @       @       @       @      �?      �?݌S���?�B����?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @-h#���?��_*>�?                                              �?       @      �?                                       @       @              �?       @m��W�?T�P{��?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @nC��x�?67�K�?                      �?      �?(�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @����[�?��[	�k�?                                �@�6�?      �?       @      �?                       @               @       @              �?       @��¯�D�?�B#X�h�?              �?                 �
���?      �?              �?                                       @       @              �?       @�`ph>�?�:B;�:�?                      �?                      �?                                                       @                              @��J�ć�?���[4q?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�%��}�?��X����?              �?      �?        ��ۥ���?      �?       @      �?       @                                               @      �?      �?�AQ�s��?`X���?      �?                        �ԓ�ۥ�?      �?                       @       @       @                              �?              @q���Y�?������?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�X����?̜�#��?      �?              �?        �z2~���?      �?       @      �?       @               @                                      �?      @�>�MF�?�bM�J�?                      �?        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                        m+�oM�?B���Rbo?      �?              �?        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              @]����`�?�W�� �?                                ��ۥ���?      �?       @                       @               @               @      �?      �?      @���S��?���i�?                                ?���@��?      �?              �?                                                              �?       @'#��~��?�0��|�?      �?              �?      �?      �?              �?               @               @       @       @               @              @q
Sb���?�kh����?      �?              �?        ��ۥ���?              �?                       @                       @       @       @               @*L����?��J�i��?      �?              �?        (�K=�?      �?       @      �?       @       @       @       @       @       @       @              �?(��E��?X�@�_�?      �?                        �K=��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����'t�?�=JUc�?      �?                        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?        ^��Z��?T�P{��?      �?                        �z2~���?      �?       @      �?               @                       @       @              �?      �?#s�g�L�?����n�?                      �?      �?6���?              �?               @               @       @       @       @       @              @<�RG�m�?��Ǝ���?      �?      �?      �?        3~�ԓ��?      �?              �?                                               @              �?      �?������?�{+��2�?                      �?      �?6��9�?      �?                       @       @                       @       @      �?                ��8j��?���3�?      �?              �?              �?      �?       @                       @       @               @       @       @                :�X�?�p��%J�?              �?                ��RO�o�?      �?       @      �?                                                              �?       @j�����?"�N#Կ?      �?                      �? �
���?              �?                       @                       @              �?      �?        '���G��?�KI�ܯ�?      �?              �?        ��Vؼ?      �?       @      �?       @                                       @              �?       @��r�9�?�����?              �?                3~�ԓ��?      �?       @      �?                       @                       @              �?        �=����?P��Bb�?                                6��9�?              �?               @       @       @                                                �^!ї�?q�w@o�?                      �?      �?�ԓ�ۥ�?      �?       @      �?       @       @       @       @       @       @       @              �?)��|�?�?������?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @����[�?k�7�O�?      �?                        ��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?�+��ޒ?                              �?�'�K=�?      �?              �?               @                               @              �?        >�� Q��?gw'tZy�?                      �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?�F�'1��?                                ���V،?      �?       @      �?                                               @              �?       @1v�z�?-�.ٴב?                                �'�K=�?      �?       @      �?                                                              �?       @�J���?�v_�)�?      �?      �?                �RO�o��?      �?       @               @       @                               @      �?      �?       @�{'Y��?g�r��?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                       @1[�yj�?k���>[�?      �?      �?      �?        ���V؜?      �?       @      �?               @       @               @       @              �?       @r@����?A}u�/��?      �?                        ��V��?      �?       @                       @                                              �?        �5A .�?��T dQ�?                                ���V؜?      �?       @                                                                      �?      @�{B���?B;�m,P�?                      �?      �?!�
���?      �?               @      �?      �?      �?      �?      �?      �?       @              @8�]�FR�?�Z���ս?      �?                                      �?              �?                                                              �?       @X-�r�?�3�
'x?      �?                        6��9�?      �?              �?                                       @       @              �?       @���¯�?�36��?              �?                              �?              �?                                                              �?       @'#��~��?KnJEx?      �?              �?      �?F���@��?      �?              �?                                                              �?        ��j1v�?�/��C,�?      �?              �?        {2~�ԓ�?      �?       @      �?               @                       @       @              �?       @��G��q�?�BAM�<�?      �?                                      �?       @      �?                                                              �?       @�ae��	�?��	�z?              �?                ��.�d��?      �?       @               @               @                               @                G�%��}�?���{��?              �?                              �?              �?                                                              �?       @�l	�Y�?�-˽x?      �?              �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�d�Q�ϐ?׿����?                                ���V،?      �?       @      �?                                       @       @              �?       @4�돗��??3�z�n�?      �?              �?        v�'�K�?      �?       @                                       @               @                       @<�$0�	�?��<�#[�?                      �?        ���V،?      �?              �?                                                              �?       @3NaJ̖�?������?      �?              �?      �?6��9�?              �?               @       @                                              �?      @H*��E�?o9#{kx�?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?                      @�%��}�?����?      �?                        ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      @��1�~?���h|?                      �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?                        �U�����?���	�Ѳ?      �?              �?      �?��ۥ���?      �?       @               @       @               @                      �?      �?      �?���J��?\?N�0w�?                              �?[as �
�?      �?       @      �?                                       @                      �?      �?&�1�L��?��I	.��?      �?      �?      �?        ܥ���.�?      �?       @      �?                       @                       @              �?      �?�5A .�?f=4���?      �?                        6��9�?              �?                                                                      �?        qi��|��?����`��?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?              �?       @�^W-��?%�eXg�?              �?      �?              �?      �?       @      �?               @       @               @       @      �?              �?e0
84��?SW����?      �?                        �ԓ�ۥ�?      �?       @      �?       @       @       @       @                              �?      @��C���?������?      �?                        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�^W-��?G�Zlno?      �?              �?        ܥ���.�?      �?       @                       @       @                       @      �?      �?      �?@y4���?]@G�?      �?      �?      �?        ��RO�o�?      �?              �?                                                              �?       @@y4���?>hJ7o�?      �?                        �ԓ�ۥ�?      �?                       @               @       @       @                      �?       @l?C؋��?d�,���?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @�፿Po�?��߄3�s?      �?                        �@�6�?      �?                                       @               @       @              �?       @�vAIE�?���e*|�?      �?                        �ԓ�ۥ�?      �?       @      �?       @       @       @               @       @       @      �?      �?b/��:�?U�Oˊ^�?      �?      �?                p�z2~��?      �?              �?                                                                      �?�¯�Dz�?�I?�>P�?                              �?�@�6�?      �?                       @               @                       @      �?              @�\d����?��9գw�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?1[�yj�?�ݏљ?                                ?���@��?      �?                       @                                                      �?        �Po���?�h�b���?                      �?      �?�
��V�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?g�)L�ٲ?���<9�?                      �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @                �'�F7�?UKқ]N�?      �?              �?      �?�K=��?      �?       @      �?                       @                       @              �?      �?�^!ї��?.�����?      �?                                      �?                                       @                                      �?      @O�)���?��.��)m?      �?      �?                �'�K=�?      �?       @      �?                       @               @       @              �?       @S}䛌8�?�֌�z��?      �?              �?      �?      �?      �?       @               @       @       @       @                       @              �?���q%�?��e*|t�?                      �?      �?      �?      �?       @                       @               @       @       @       @      �?       @L���S�?+�ل��?                                3~�ԓ��?      �?                                       @                       @      �?              �?��l	��?P-�2��?                                              �?                                                                                      �?�7�B�]�?#��=�g?              �?                ���V؜?      �?       @      �?               @                                              �?       @)�tN|x�?Ř�>�?      �?              �?      �?�'�K=�?      �?              �?       @                                                              @��8j��?��+��?                      �?      �?	��V��?      �?              �?       @                       @       @                               @�፿Po�?����>��?                                ?���@��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�p�Ȭ?K���M��?      �?              �?        ���V؜?              �?                                       @                              �?       @�\d����?daL��[�?      �?              �?        ���V،?      �?                               @               @               @              �?      @�ć7�B�?TS�[Z��?      �?      �?      �?        P�o�z2�?              �?               @       @       @                               @      �?       @��a/�?-�2���?      �?                        �'�K=�?      �?       @      �?                               @       @               @      �?      �?��ǰ2��?6�C��=�?                      �?        ��RO�o�?      �?       @      �?                       @                       @                        �
����?>�M'��?      �?      �?      �?        ��RO�o�?      �?       @      �?               @       @               @       @              �?       @���vA�?�Ȱ/�?                      �?        ���V،?      �?              �?                                                              �?       @���S��?���A��?                      �?        (�K=�?      �?       @               @               @       @                       @              �?o��R��?
�`����?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @�Y;���?�E&��3�?      �?      �?                $Zas �?      �?                       @                       @                      �?              @�d�#��?F��s���?      �?              �?      �?�6��?      �?       @      �?                       @       @       @               @      �?        p2��g�?���1]��?      �?              �?      �?{2~�ԓ�?      �?              �?                       @               @              �?      �?       @H*��E�?��z����?                                �]�����?      �?       @      �?       @       @       @       @       @       @       @              �?�c=kg��?8B�X��?      �?      �?      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                3�$0�	�?e9F){��?      �?      �?      �?        �K=��?      �?       @      �?                                       @       @              �?      �?�<݌S�?/��i�`�?      �?              �?        �
��V�?      �?                       @       @               @                                      @I8O�)�?�F}��?                      �?      �?p�z2~��?      �?       @               @       @                       @       @      �?               @��T�&�?�C����?                      �?        >�]���?      �?       @      �?       @       @       @               @       @      �?                �9ֳv&�?M좤�}�?      �?              �?        �K=��?      �?              �?       @       @                               @      �?      �?      �?���l	�?��>� K�?                                ���V؜?      �?              �?                       @       @                                      �?���U���?c,kR!|�?      �?              �?        (�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                qi��|��?T=��c�?                      �?      �?ܥ���.�?      �?       @                       @               @       @       @       @               @��<݌�?g\�8�q�?      �?                        ���V،?              �?                                                                      �?       @?�]�FR�?>����q?      �?              �?      �?[as �
�?      �?       @                                                       @                        �3i�ae�?'��넯�?      �?                        ��.�d��?      �?                       @       @                       @               @      �?      �?�1���?-GB���?                      �?      �?�K=��?              �?                       @       @       @       @       @       @      �?       @!s�g�L�?PoS�Q+�?                                {2~�ԓ�?      �?       @                               @       @       @       @      �?      �?      @�F���?*�-����?                      �?        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @                ���'tX?7J�����?      �?                        ���V؜?      �?              �?                                                              �?      @p�l�?���Wҗ?                                �z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�r@��?/2�]��?              �?      �?        ��RO�o�?      �?       @                       @       @       @       @       @                       @�'�F7��?ֵ#��?      �?      �?      �?        Zas �
�?      �?       @      �?                       @               @       @              �?       @ /�Q���?M���+�?      �?                      �?                      �?                                                                              @)���O�?�+;p&kD?                      �?      �?�ԓ�ۥ�?      �?                                       @       @                      �?      �?      �? J�hY�?���yӷ�?      �?                        ���V؜?      �?       @      �?                                                                      @�N���?��_%�|�?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?      �?W����?<V��T��?      �?              �?        �]�����?      �?              �?                       @               @       @              �?      �?c9�W�?h=�K��?      �?                        	��V��?      �?                       @       @                                              �?      �?�#�6���?��.�D
�?                                �@�6�?      �?                                               @                              �?        O�)���?�ؐ^�?      �?              �?      �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�U����|?��iiǔ�?                                {2~�ԓ�?      �?       @      �?                       @       @       @       @      �?      �?      �?�<5���?V7����?                      �?      �?[as �
�?      �?       @      �?               @                               @              �?       @F�*�A6�?�Mܬ��?                                ��RO�o�?      �?              �?       @       @       @       @               @       @              @�۴���?i��l���?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?       @               @       @       @       @      �?      �?      @�.�c�?�l��?      �?      �?                ��.�d��?              �?                       @                       @       @              �?       @���w��?gte�4��?                      �?      �?��ۥ���?      �?                       @                                                              �?�'�F7��?���ч�?                                ��ۥ���?      �?                       @       @       @       @       @       @      �?                z�Τ=��?J�!9�
�?      �?              �?        ��Vؼ?              �?                                                              �?                ò
n�ͭ?��3.z�?                                ��Vؼ?              �?                       @                               @                       @�1���?}���?                      �?        �ԓ�ۥ�?      �?       @      �?                       @       @       @       @       @                �������?��lת�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @F��1��?��1�SH�?                                ��Vؼ?      �?              �?                                       @       @              �?      @Z;��V�?ٮS����?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                       @����'t�?�>�!�+?              �?                �@�6�?      �?       @               @                                                      �?       @�N�����?*|����?      �?              �?        �K=��?      �?       @      �?               @                       @              �?      �?        Z;��V�?"�b�aW�?              �?      �?        �ԓ�ۥ�?      �?              �?       @       @                               @      �?              �?�Ήo��? Ef��J�?                      �?        ��ۥ���?      �?       @      �?                                       @       @       @      �?        %0�	�?\b��a?�?      �?              �?      �?�K=��?      �?              �?                                       @                               @c=kg��?�)@���?      �?                      �?��RO�o�?      �?                       @       @               @                      �?              �?�����f�?G�nc�?      �?              �?        �'�K=�?      �?       @      �?                                               @              �?        o��4�u�?�J[���?              �?                ��Vؼ?      �?       @      �?                                                              �?       @9ֳv&��?(�Orvر?                      �?        �o�z2~�?      �?              �?       @               @       @       @       @      �?      �?       @��0%f�?h��z"Z�?              �?                ���.�d�?      �?       @      �?       @               @       @       @       @              �?        ��-��?�����0�?              �?                e�v�'��?      �?       @      �?               @                                              �?       @�?^���?6��p�?                      �?      �?�'�K=�?      �?       @               @               @       @       @       @       @      �?       @�s��2�?w����?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?M:'>��?r�@�f�?      �?                        ���V،?      �?              �?               @                                              �?       @F��s��?���c�ƍ?                                F���@��?              �?                                                                                ?�]�FR�?���<9�?                      �?      �?p�z2~��?              �?               @       @       @               @       @       @      �?      �?ٴ��I��?6���N�?                      �?        p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�.h#��?.B��2�?                                �'�K=�?      �?              �?                                       @                      �?       @��䶺O�?A�n{�w�?                                �ԓ�ۥ�?      �?       @      �?                               @               @              �?       @C)-���?�����?      �?                      �?�'�K=�?              �?               @       @       @       @                              �?      @�{'Y��?�f���?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @              �?+�oM��?�}�i�V�?                                              �?              �?                               @       @       @              �?       @�>|]��?7��{5�?      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?       @                m+�oM�?��U���?                                ?���@��?              �?                                                                      �?       @h#���?���b��?      �?      �?                H���@��?      �?       @      �?                                       @       @              �?       @Aʾ����?�]�hZ�?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                        ����[�?H���e�?      �?                        6��9�?      �?       @      �?                               @       @       @                        ��w�ӥ�?�g[��?      �?      �?                �K=��?      �?       @               @       @               @                       @      �?        ���>|�?(_��?�?                                ���@��?      �?       @      �?       @       @               @       @       @       @      �?       @H���<�?>��m�?      �?      �?      �?        ���.�d�?      �?       @      �?                       @       @       @       @       @               @1@�bѲ�?=$�@�?      �?                        F���@��?      �?              �?                       @                                              @�k�.M��?("���?      �?                        �V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����[�?�\.�E�?                      �?      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @�U�����?nS�<��s?      �?              �?      �?�RO�o��?      �?       @      �?               @               @       @       @              �?        Wc"=P9�?Q�Ő���?                      �?      �?�z2~���?              �?               @                               @       @              �?        jg����?�@����?      �?              �?      �?p�z2~��?      �?       @               @               @       @       @       @      �?      �?      @y4��0�?�y�ek�?      �?                        F���@��?      �?       @      �?                       @               @                      �?      �?�G�Ɉ��?�_5{%�?                      �?        P�o�z2�?      �?       @               @                       @                      �?                �C��x�?��V�8�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?��n�X�%?              �?      �?        ?���@��?      �?       @      �?       @                               @       @              �?       @��l	��?ʑ�m�?                                ���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @,1[�yj�?4�y���?                      �?      �?(�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?        ���O��?a��j�s�?              �?                              �?       @                                                                              @�Po���?&��=mn?      �?                        �V�H�?              �?               @                                              �?      �?        _ph>׿?���lF��?                                              �?              �?       @                               @       @              �?       @IE����?;}m[&�?      �?      �?      �?        F���@��?      �?              �?               @               @               @              �?        B����?�IZ�y��?                              �?(�K=�?      �?       @               @       @               @                       @               @��`ph�?���'.��?                                �'�K=�?      �?       @               @       @       @                                      �?        ��@���?,t];`�?      �?              �?        �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?Rp�l?c} �?      �?                        �'�K=�?              �?                               @       @       @       @       @              �?�R,Z�?,��҆��?      �?              �?      �?���V؜?      �?                                       @                                      �?       @��"X~P�?$K�^˥�?                                ?���@��?      �?       @      �?               @                                              �?      @������?�ׅ!�?                                              �?              �?                                                                        K��a�?��]�x?      �?      �?      �?        ���@��?      �?       @      �?       @               @               @       @       @      �?      �?)���G��?�ˍ ��?                                	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @����[�?���Վȣ?      �?              �?        ?���@��?      �?       @                               @               @                               @�U:'�?>�9�T�?      �?                      �?�K=��?      �?       @      �?       @       @                       @       @      �?      �?       @.�c=�?]�`~�?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?              �?       @��N�ԑ?wm��П?              �?                �o�z2~�?      �?       @      �?                                       @              �?               @#���?xc^L!>�?              �?      �?        �'�K=�?      �?       @      �?               @       @                       @                      �?��1��?=�~ʯ�?      �?              �?        ���V،?      �?       @      �?                       @               @                      �?       @؋�ߵN�?T��S�	�?                                6��9�?      �?       @      �?       @                               @       @              �?       @]d�����?�����1�?      �?                        ��ۥ���?      �?                       @               @       @       @       @              �?      �?��.h�?&hR���?      �?              �?      �?���Vج?      �?               @      �?      �?      �?      �?      �?      �?      �?              @Y�)L�ْ?i
�69V?      �?      �?      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �d�Q�ϰ?�uy9 ��?      �?      �?      �?        !�
���?      �?       @      �?       @               @                       @      �?      �?        be��	�?(7D����?                                �V�H�?      �?              �?       @       @       @               @              �?      �?      �?�:��?(�:P'�?      �?              �?      �?      �?              �?               @       @       @       @       @       @       @      �?        ��a/�?�����'�?                      �?         �
���?      �?              �?                               @               @                      �?>�� Q��?��l��?              �?                ���V،?      �?              �?               @                       @                      �?        :]��#��?�I�.�?      �?              �?        �]�����?      �?                       @                       @                      �?      �?      �?��s��2�?��q���?      �?                        ��ۥ���?      �?       @      �?                                               @              �?       @�iŽ�,�?�whc�?              �?                �'�K=�?              �?                       @       @               @       @              �?       @jL�*g�? �1���?                      �?        >�]���?      �?       @      �?               @       @       @                                       @ J�hY�?������?                      �?        �'�K=�?      �?       @      �?                                               @              �?       @ ʣ��8�?�����
�?                      �?        {2~�ԓ�?      �?       @      �?                               @                              �?      �?���Z�K�?�
����?              �?      �?      �?>�]���?      �?                       @                       @       @       @       @      �?      �?�ht3N�?�:o[�?              �?                F���@��?      �?                               @       @                                      �?       @R��'�F�?�8[�:�?                      �?                      �?              �?                                                              �?       @� �;�$�?w�ו�w?                                �'�K=�?      �?              �?                                       @                      �?        M+�d��?`�y�Q�?      �?      �?      �?        �]�����?      �?              �?                                       @       @              �?        �d�#��?�`O\�?      �?      �?                ���V؜?      �?              �?                                       @                      �?       @ȕ�=��?�=�t��?                                              �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?J���q'?                              �?�ԓ�ۥ�?              �?                                                       @              �?       @SUUUUU�?������?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?                      @����[�? �<$3?                      �?      �?3~�ԓ��?      �?                       @       @       @       @               @       @              @�Ɉ����?Z������?      �?      �?      �?        �@�6�?      �?       @      �?                       @               @       @              �?       @!ї�V��?��LmQ�?              �?      �?        (�K=�?      �?       @      �?               @               @       @       @      �?      �?        ��+	��?�Ö���?      �?                        ���Vج?      �?                                       @               @       @              �?       @���"X~�?��b�Z�?      �?                        $Zas �?              �?                                       @               @              �?       @�*�A6w�?C�#����?      �?              �?      �?�
��V�?      �?       @      �?                                       @       @      �?                Gm?C؋�?$a����?                      �?      �?�'�K=�?      �?              �?                                       @       @              �?      �?4��0%�? ��'9�?                      �?        ���V؜?      �?       @      �?               @                               @              �?      �?�V�;�R�?&��y|�?                                �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                        �፿Po�?4|����?                                !�
���?      �?              �?                                       @       @      �?              �?d�Q���?A��Ou�?                                �'�K=�?      �?                       @                                                      �?       @h#���?� )2�|�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?�^/��"?      �?              �?      �?H���@��?              �?                       @                       @       @      �?      �?        ��>|]�?��2(���?                                �'�K=�?      �?       @               @                       @               @                       @f��	��?c[�c�?              �?                [as �
�?      �?       @      �?               @                       @       @              �?       @k1v��?��,�(e�?      �?              �?        (�K=�?      �?       @      �?               @       @       @               @       @      �?        ]d�����?���i�A�?                      �?      �?              �?              �?                                       @                      �?      @���w��?�N�-�|?      �?                        	��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�m��W�?�J��H.�?      �?              �?        (�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?m+�oM�? *��j��?      �?                      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @m+�oM�?���4��?                      �?         �
���?      �?                               @       @       @       @       @                        EDDDDD�?S"G�Zl�?                      �?      �?��.�d��?      �?       @      �?                       @               @       @      �?                ;�RG�m�?$X�h`��?      �?              �?      �?�6��?      �?               @      �?      �?      �?      �?      �?      �?                       @�X����?g�[��?      �?              �?        �K=��?      �?       @      �?               @       @                       @       @      �?       @�yjH��?`5{%r�?                      �?      �?�D+l$�?      �?                               @       @       @       @       @       @                �:]���?㇔&�[�?              �?                 �
���?      �?       @      �?       @       @                               @              �?       @���`p�?�)�M�?                      �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?      �?                �%��}�?7�O�k�?                                �K=��?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?��]Q�T�?      �?                        p�z2~��?      �?              �?               @       @                       @              �?       @�r�9ֳ�?��6d�?      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?-h#���?�����?      �?      �?      �?        v�'�K�?      �?       @      �?                               @       @       @              �?      �?��_���?ŵIbBN�?                                �ԓ�ۥ�?      �?              �?       @                                                      �?       @/M��o2�?��:��?                      �?      �?��.�d��?      �?       @      �?               @       @               @              �?      �?      �?��.h#��?�)SB3N�?                      �?      �?ܥ���.�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�%��}�?�F}���?      �?      �?      �?              �?              �?               @       @       @       @       @       @       @      �?        ^�ti���?>�к~;�?      �?                        $Zas �?      �?       @                       @               @       @              �?      �?       @+�oM�?4C�Lޣ�?      �?              �?        p�z2~��?      �?       @      �?               @                                      �?      �?       @��䶺O�?)�p���?      �?      �?                P�o�z2�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?��N�ԑ?Ƌ��|W�?      �?                        !�
���?      �?       @      �?               @                                                        �����?Q(,	�?                              �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?              �?       @�፿Po�?q����?      �?              �?      �?�V�H�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        #w\I`ޓ?8Wꈝl�?      �?                        �'�K=�?      �?                                                               @              �?      �?�`ph>�?�ЄŨ?                                p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @              @����[�?kA`n�Y�?      �?      �?                              �?              �?                                                              �?       @�=�� �?m[����x?                                SO�o�z�?      �?              �?               @       @       @       @       @              �?        .�c=�?�z����?              �?      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?        �8j���?VU�%7��?      �?                         �
���?      �?       @      �?       @       @                       @                      �?      �?T��%��?|9�=7�?                      �?        3~�ԓ��?      �?       @      �?               @       @       @       @       @       @      �?        /�Q����?��Ntm1�?                                ���Vج?      �?              �?                               @                              �?      @�B�]�F�?����F}�?      �?              �?        ,l$Za�?      �?              �?                                       @       @      �?      �?        �ߚ ��?�o�$6�?                      �?      �?v�'�K�?      �?       @      �?       @       @       @               @       @       @                /�Q����?��W�?                                p�z2~��?      �?                                       @                                      �?      �?���!���?b[�c��?                                              �?                                               @                              �?       @��̱��?t!��o?                      �?        ��V��?      �?               @      �?      �?      �?      �?      �?      �?       @                ,1[�yj�?�>0�7�?      �?              �?      �?�'�K=�?      �?              �?                       @               @       @              �?       @&���[�?8�R��?                                ���V؜?      �?                                       @               @                               @(-���?0/�ې?      �?              �?        ��ۥ���?      �?       @      �?       @       @       @               @               @      �?       @�$K!��?{�1�?��?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?                       @               @       @              �?      �?�E�X���?H��x���?                                ���V؜?      �?              �?                                       @                      �?       @�~5&��?��m�;�?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?����[�?�����ww?      �?      �?                �'�K=�?      �?              �?                                               @              �?       @)�tN|x�?<v��_��?                                [as �
�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�X����?	^��ڠ�?                                              �?       @                                                                      �?        uN|x�/�?�Lhe:rm?                                Zas �
�?      �?       @      �?       @       @       @       @       @       @      �?      �?       @��!����?��$�!�?      �?                        �'�K=�?              �?                       @               @                                       @���7q�?��, �?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�j1v�?���5�.�?                      �?      �?[as �
�?      �?                       @               @       @       @       @      �?      �?      @�b��!�?���"x��?                                �D+l$�?      �?       @      �?               @                       @       @              �?       @:'>���?�xP���?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        ��^<��?��E I�?      �?                        p�z2~��?      �?              �?                                       @       @              �?       @����?�d�?      �?              �?      �?�K=��?      �?       @      �?       @                       @       @       @       @                M�cX�~�?NZ[�?                                �D+l$�?      �?       @               @       @       @       @               @      �?              �?��*��?�Y����?                              �?�@�6�?      �?                                                                                        ���8�)�?��W����?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @                s����?C�.ٴ��?                      �?      �?(�K=�?      �?       @               @       @                       @               @      �?      �?�c9�?�)���?      �?                        H���@��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @nC��x�?�Jte�?      �?              �?      �?H���@��?      �?              �?                               @       @                               @>�� Q��?(�����?      �?                      �?{2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ���C�?�?�)�?      �?              �?      �?�]�����?      �?              �?       @                                                                �N���?7l��Z��?      �?      �?                              �?       @      �?                                                              �?       @�6��`��?5� ��kz?      �?      �?      �?        �ԓ�ۥ�?      �?       @      �?               @       @                       @              �?        KS}䛌�?��'�?              �?      �?        v�'�K�?      �?       @      �?               @       @               @       @      �?              �?M�cX�~�?L����?      �?              �?        �
��V�?      �?                       @       @       @                               @               @,ZV���?�w���?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �??�]�FR�?�f��e�?                                	��V��?      �?              �?                                                              �?       @�¯�Dz�?M�G5���?              �?                ���.�d�?      �?       @                       @       @       @               @                      �?�k�.M��?����=��?      �?      �?                ���@��?      �?       @               @       @                       @                      �?        3NaJ̖�?��[W�_�?      �?                        SO�o�z�?      �?       @      �?               @                       @       @              �?       @۴��I��?�?.��k�?      �?                        ��Vؼ?      �?                                                                                      @�=�� �?���-wZ�?              �?                �D+l$�?      �?       @      �?       @       @       @                                      �?       @�d�#��?
z��w:�?      �?              �?      �?p�z2~��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @)���O�?�O,�o�?      �?                        ��RO�o�?      �?              �?                                       @       @              �?       @�J���?��z�?      �?              �?      �?,l$Za�?      �?                               @       @       @                              �?      @��+	��?�A��t�?      �?                        6��9�?      �?                                               @       @                      �?      �?�+$���?B�:���?      �?              �?        ���.�d�?      �?              �?       @       @               @       @       @       @      �?      �?�#�d�Q�?8�sLzR�?      �?                        ��ۥ���?      �?       @      �?       @       @       @       @       @       @      �?      �?        �0%fK8�?p�]F��?                      �?        ��RO�o�?      �?       @      �?               @                       @       @              �?      �?ʣ��8��?�l���?                                F���@��?      �?              �?                                       @                      �?      @������?�����?              �?                              �?       @      �?                                                              �?      @�@ʾ���?�����Mz?                      �?        �V�H�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        h#���?�/HC��?                      �?        �K=��?      �?       @      �?                                       @       @              �?       @[�yjH�?�RH���?                      �?      �?      �?      �?       @                               @               @       @       @      �?        �z�����?"���?                      �?      �?���@��?      �?               @      �?      �?      �?      �?      �?      �?       @                ����[�? �°�?      �?              �?        �V�H�?      �?               @      �?      �?      �?      �?      �?      �?                       @�X����?Y���?      �?      �?      �?      �?�]�����?              �?               @                                       @                      @=Q�s���?W�~Fr�?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @               @      �?      �?)����?6�8���?      �?                        ��Vؼ?      �?       @      �?                                       @                      �?       @��>|]�?7V$�ڵ?      �?                        SO�o�z�?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�%��}�?�s�=�?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?      �?              @8�]�FR�?�w���Qk?      �?              �?      �?�K=��?      �?       @      �?               @       @       @       @       @       @      �?        �f���?��̩��?      �?                        ?���@��?              �?                               @                                      �?       @3�$0�	�?�ͺ�ʏ�?      �?                      �?              �?                                                                              �?       @?y4���?_�<$3h?      �?      �?      �?        6��9�?      �?              �?       @                                                               @���H*�?�	r-��?      �?      �?                3~�ԓ��?      �?       @      �?                       @                                      �?      �?����?F-�m4�?                                SO�o�z�?      �?                       @               @                                              �?�
n���?7gA����?      �?                      �?�]�����?      �?       @      �?               @                       @                      �?      �?R��'��?\�J���?      �?                        �ԓ�ۥ�?      �?       @                               @       @       @       @      �?      �?      �?��-�jL�?��6���?      �?                        ?���@��?      �?                                               @       @                      �?       @|䛌8j�?8�^�?�?      �?      �?      �?                      �?       @      �?                                                              �?       @�u�b���?P��,�Gz?                      �?      �?{2~�ԓ�?      �?       @      �?               @       @               @                      �?      �?�*���?$j���?      �?                         �
���?      �?       @      �?                                               @              �?       @��x�]��?z�/HC��?      �?                        �'�K=�?              �?               @               @               @       @              �?       @N��b��?8��"�v�?      �?      �?      �?        ��.�d��?      �?       @      �?               @       @               @       @      �?      �?        ����Z��?���Վ��?      �?                      �?���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?�J�Tt�r?                                �z2~���?      �?              �?       @       @                       @       @      �?      �?       @��'t �?�M���|�?                                �@�6�?      �?                       @       @                                                       @��s��2�?V%$��?      �?                        ��V��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�%��}�?y>���?              �?                ���V؜?      �?              �?                                                              �?       @p�l�?U�����?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @      �?        8�፿P�?�����?                      �?        ��V��?      �?       @      �?               @       @       @       @       @       @      �?        �*�A6w�?:̫�?              �?                ��.�d��?              �?                       @       @       @       @                      �?       @9��_���?_��=R��?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?��;�N�?                                ���Vج?      �?               @      �?      �?      �?      �?      �?      �?              �?      @���@��?��_�4�?      �?                        ?���@��?      �?              �?                                       @       @              �?       @�R,Z�?�Q&5�ɤ?      �?                        �@�6�?      �?                               @       @       @                              �?       @I8O�)�?���Վȳ?                                ��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��+$��?��%ٷ?                      �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        Y�)L�ْ?7t��(��?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?.-˽h?      �?                        ���.�d�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�%��}�?�o�/
�?                      �?      �?��ۥ���?              �?               @       @               @       @       @       @              @��?y4��?B���~y�?      �?              �?        F���@��?      �?       @               @                                       @              �?       @3���O�?����?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?b:���9[?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @�'�F7�?O���&?      �?                        p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?       @                1[�yj�?U��"2M�?      �?              �?        p�z2~��?      �?       @      �?               @       @       @       @       @              �?       @�C��?Y�r�{��?      �?              �?      �?(�K=�?              �?               @               @       @       @       @       @                ��¯�D�?!���x�?                                �D+l$�?      �?       @               @               @               @       @      �?      �?      �?���Up�?�e{&��?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?               @                       @                      �?        h{����?7D���5�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @8�]�FR�?����d!?                      �?      �?6��9�?      �?                                       @                                      �?        �7q���?�~K+��?      �?      �?                ܥ���.�?      �?       @      �?               @                       @       @      �?      �?       @�$K!��?���1s�?      �?              �?        SO�o�z�?      �?       @      �?               @       @               @                      �?        Ž�,u��?]1��?                                �ԓ�ۥ�?      �?       @               @               @                                      �?      @%��}��?�6�Q��?      �?                        �@�6�?      �?                       @       @                                              �?        �yjH��?/��O��?                                �@�6�?      �?       @      �?               @                       @       @              �?      �?䛌8j��?J���+'�?      �?      �?      �?        �'�K=�?      �?       @      �?                                               @              �?       @�H*���?',	F�?      �?              �?        ���Vج?      �?       @      �?               @               @                              �?       @��3i�a�?Dl�{;��?      �?      �?      �?      �?���@��?      �?       @               @       @       @                       @       @      �?        _W-��?�r5�?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�U�����?P���?      �?              �?      �?�@�6�?      �?                       @                                                      �?       @���w��?ٖ �P[�?                      �?        �z2~���?      �?       @      �?                       @                       @                      @�
����?�#�~N��?                      �?      �?,l$Za�?      �?               @      �?      �?      �?      �?      �?      �?                      @�X����?�|1$i~�?      �?              �?      �?�'�K=�?      �?       @                               @       @                              �?        .��:]�?��K#5�?      �?              �?        Zas �
�?      �?       @      �?               @       @               @       @              �?       @��+	��?W�� �?      �?              �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @nC��x�?-�2�ý?      �?              �?      �?P�o�z2�?      �?              �?       @       @               @               @       @                {]�;x�?*����?                      �?        ��V��?      �?                       @               @       @                       @              �?R�����?ۅ�{�X�?      �?              �?        �o�z2~�?              �?                                       @       @               @      �?        <�RG�m�?�����?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�U�����?FPeB�?      �?                      �?Zas �
�?      �?       @               @       @                               @              �?       @%�yO�0�?1�!�:u�?                      �?      �?�@�6�?      �?       @      �?               @       @               @                      �?      @z����"�?!�Z𫉭?      �?              �?        �'�K=�?      �?       @      �?               @                                              �?        ��̱���?�'Tn'��?      �?              �?      �?!�
���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�፿Po�?�, =�?                                ��V��?              �?               @               @       @       @       @       @              �?V�&#��?� 0���?      �?                        �ԓ�ۥ�?      �?       @      �?               @               @       @       @      �?      �?        s[ݧ���?mRI4�?              �?      �?        �]�����?      �?       @      �?                       @       @       @       @      �?      �?       @E�Ήo�?q֜�#��?                      �?      �?��RO�o�?      �?       @      �?                               @       @                      �?       @嶺O_�?u�m�E��?      �?              �?      �?�D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?E�(Ţe�?y�\�V�?                                ���@��?      �?              �?                       @       @               @       @      �?        +�oM��?�����?      �?              �?      �?,l$Za�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @��+$��?f����?      �?                        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                      @F��1��?v[�ɎL�?      �?              �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              @����'t�?r��� �?                                ?���@��?              �?               @               @       @               @                      @�rv��?uD{@O��?      �?              �?      �?H���@��?      �?       @      �?               @       @               @              �?      �?       @be��	�?]��O$��?      �?      �?                ��Vؼ?      �?       @      �?               @                       @       @              �?      �?�E�X���?	������?                              �?���V،?      �?               @      �?      �?      �?      �?      �?      �?      �?                ���@��?����bb?                                ��Vؼ?      �?              �?                                                                       @������?7
��O�?                      �?        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����'t�?�b�.O�?      �?                      �?���V؜?      �?                       @               @                                              @������?pg��%e�?                      �?      �?6��9�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @Rp�l?����ј�?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @m+�oM�?����b�?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����`�?���V�x?      �?              �?      �?�
��V�?      �?              �?               @       @       @       @              �?                �J���?�A@�QN�?      �?                        �]�����?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @��N�Ա?%�|�-�?      �?                      �?              �?                                                                                       @����e�?���W�g?                      �?      �?	��V��?      �?       @       @      �?      �?      �?      �?      �?      �?                      @ò
n�ͭ?�9�T�?              �?                �ԓ�ۥ�?      �?       @      �?               @               @       @       @              �?      �?D)-�?����g�?      �?              �?      �?�
��V�?      �?                                       @       @                       @      �?      �?
84���?�����?                      �?      �?�
��V�?      �?                       @       @                                                       @�yjH��?{��u��?      �?                        F���@��?      �?                                                                              �?        �d�Q���?�h�/k�?      �?              �?      �?3~�ԓ��?      �?              �?                                                              �?        ����e�?|^D�i3�?              �?                6��9�?              �?                                       @                              �?       @3�$0�	�?�}M"	�?              �?      �?        SO�o�z�?      �?       @      �?               @       @               @                      �?       @X~PT��?"��$���?      �?      �?                ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                        n��W�?t����΁?      �?                        ��.�d��?              �?               @       @       @       @       @       @       @              �?�C��?��#K�}�?      �?      �?      �?        F���@��?      �?       @               @       @               @                                       @�ć7�B�?�����?                      �?        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?                        �፿Po�?Hzb�?      �?              �?        ��RO�o�?      �?       @      �?               @               @               @      �?                �Wc"=P�?�O4���?      �?              �?      �?��RO�o�?      �?       @               @               @       @       @       @                       @1v�z�?2�r����?                      �?        �D+l$�?      �?       @      �?               @               @       @                      �?      �?=���&�?ق�����?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?                        nC��x�?��NIDM�?      �?                        ?���@��?      �?                                               @                              �?      @]<��u��?0x�rҮ�?                                              �?              �?               @               @       @                               @����c�?��nh:�?      �?                                      �?       @                                                                              @ئ�N��?X2��3n?      �?                        ?���@��?      �?       @                                                                              @+���?y�?<ޣT�0�?                      �?      �?p�z2~��?      �?       @               @               @               @       @       @              �?��'�F7�?��}��?                      �?      �?��V��?      �?       @      �?       @       @               @       @               @      �?      �?��?y4��?H�����?                                6��9�?      �?       @      �?                               @       @       @                      �?��'t �?��#��?      �?              �?      �?�@�6�?      �?                       @       @       @                              �?      �?        �5\.2��?���~Vh�?                                �ԓ�ۥ�?              �?                                                                               @�^W-��?�[ËLr�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @n��W�?�^/��"?                                ���.�d�?      �?       @      �?               @       @       @       @       @       @      �?      �?=P9��_�?����?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        t+�oM�?Gv&����?                                ���V؜?      �?              �?                                                              �?        ���U�?�d����?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?                      @m+�oM�?�?Y�?                                ��ۥ���?      �?       @      �?       @       @       @       @       @       @       @              @o��z���?!��Sk�?      �?              �?      �?Zas �
�?      �?              �?               @               @       @       @      �?      �?        �n�)L��?�;�N��?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?���C�?�HY��?      �?                        6���?      �?       @      �?                       @       @       @       @      �?      �?       @�X����?N�J���?                      �?      �?�'�K=�?      �?                       @               @       @                      �?      �?      @���+$�?{�X,�
�?                      �?        ���V،?      �?              �?       @                                                      �?       @�u�b���?���:��?      �?              �?      �?���.�d�?      �?              �?       @       @                                                       @O�)���?�ʪJ���?      �?              �?      �?>�]���?      �?              �?               @       @       @                      �?      �?      @z�Τ=��?7#��ҡ�?      �?                        �'�K=�?      �?       @      �?                                                              �?       @̖p���?�I�-�Z�?      �?      �?              �?>�]���?      �?              �?       @                               @       @      �?              �?����_�?���^�?      �?              �?      �?v�'�K�?      �?       @                               @               @               @      �?        uAIE��?�a$Y���?                                ���V،?      �?              �?                                                                       @�7�B�]�?�v<#܍?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?       @7O�)��?, Q��
�?      �?      �?      �?        F���@��?      �?              �?                                       @       @              �?       @�F��?c���T�?      �?                                      �?              �?                                       @                      �?       @��r�9��?@f3­/}?      �?      �?      �?              �?      �?                       @       @       @       @       @               @                �u�b���?�*L�ù�?      �?                        �'�K=�?              �?                                                                      �?      �?��N�Ա?;�;��ʓ?                      �?      �?�D+l$�?              �?                                       @       @       @                      �?��Kn���?: �[G��?                                              �?                                                                              �?       @Z��r�?0-V�ai?                      �?        e�v�'��?      �?       @      �?       @       @       @       @       @       @      �?      �?      @���̱�?K�_{�D�?                                $Zas �?              �?               @       @               @                      �?      �?        ~(Ţe�?/,����?                      �?      �?	��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @nC��x�?b�b����?                              �?��RO�o�?      �?                                       @               @                      �?      �?�^<��u�?���Ϸ?      �?              �?        �K=��?      �?       @      �?                       @               @       @                       @#s�g�L�?�@�1��?                      �?      �?3~�ԓ��?      �?              �?               @                       @                      �?       @J̖p���?s:�P���?      �?      �?                �'�K=�?      �?       @      �?               @               @       @       @              �?        ߚ ���?��۱���?      �?              �?      �?�'�K=�?      �?                                       @       @       @       @       @              @x�ӥ�>�?v�&
�?                      �?        ��.�d��?      �?       @      �?               @       @               @                                �q%�yO�?�x�q"}�?      �?                        p�z2~��?      �?       @                                       @                      �?                9�WH�%�?�hEN �?      �?                                      �?                       @                                                      �?      @Q,?(��?����'n?      �?                        ���V؜?      �?       @      �?                                               @              �?       @ J�hY�?�Z�m�?      �?              �?      �?>�]���?      �?                       @       @       @                               @      �?        �^<��u�?�c�"e�?      �?              �?      �?(�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?E�(Ţe�?K4�MB�?      �?              �?      �?3~�ԓ��?      �?              �?       @       @       @                       @      �?              @����_�?�����?      �?              �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�0[�yjv?H,X��P�?      �?              �?        {2~�ԓ�?      �?              �?               @       @                                      �?       @M+�d��?�BQC�?                      �?        ���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        m+�oM�?Aw��M�?      �?                        ,l$Za�?      �?       @                       @       @       @       @       @      �?      �?        UUUUUU�?��c�7�?                              �?              �?       @       @      �?      �?      �?      �?      �?      �?                      @^Zq�$K�?G�O��C?      �?              �?        ��ۥ���?      �?                       @                       @                       @                ,u�ئ�?��a?���?      �?      �?                      �?      �?       @      �?       @       @       @       @       @       @       @                ��Up�l�?0������?      �?                        ���V،?      �?                                               @                              �?      �?:�X�?�}=,`�?                                �RO�o��?      �?       @      �?               @       @               @       @       @               @�oM���?�[m�Q�?                      �?      �?6��9�?      �?       @               @       @                       @              �?               @p�l�?r��v)k�?      �?                        ?���@��?      �?       @       @      �?      �?      �?      �?      �?      �?                      @��N�Ա?�x�����?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @1[�yj�?؄�3��(?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @E�(Ţe�?#md��y�?      �?                      �?���Vج?      �?                                               @                              �?        ����[�?��S�	��?              �?                ���V،?      �?                                                                                       @�7�B�]�?i
�69V?      �?              �?        ��ۥ���?      �?       @      �?               @       @       @       @       @       @      �?      �?E7����?1$i~vT�?      �?              �?      �?�@�6�?              �?                                                                      �?       @2w\I`޳?�E(�?                      �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�፿Po�?62��_�?                      �?      �?�@�6�?      �?                                               @                              �?      @d��ht�?JuPu�?                      �?        �K=��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        9�%��}�?�Y=�T�?              �?                              �?              �?                                                              �?       @�l	�Y�?�-˽x?                                ���V،?      �?              �?                       @                                      �?       @G��q
S�?ZQ�Ő?      �?              �?      �?[as �
�?      �?                                       @       @                                      @��ǰ2��?������?              �?      �?        >�]���?      �?       @      �?                       @               @       @              �?        H���<�?l�j)��?      �?              �?      �?!�
���?      �?                       @       @               @                       @              �?����?��jG���?                      �?      �?�@�6�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @)g��1�?NN�c���?      �?              �?      �?Zas �
�?      �?       @                               @       @       @       @       @      �?        �����?�)SB3N�?      �?      �?                ���V،?      �?               @      �?      �?      �?      �?      �?      �?                       @����[�?Ǘ���da?      �?              �?        Zas �
�?      �?              �?       @       @                                                        �F���?���=�?      �?              �?      �?H���@��?      �?                       @       @               @                                      �?��U�?��k` ��?      �?                        F���@��?      �?              �?               @                       @       @              �?       @��s��2�?�25�?                      �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              @�X����?*y� ��?      �?                        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                      @1[�yj�?N����?                                �'�K=�?      �?       @               @                                                      �?      @�yjH��?�*��?      �?      �?      �?        ?���@��?      �?              �?                                                              �?       @��6���?�EQ���?                      �?        ���V؜?      �?                                                                              �?      @U:'>��?&kZ�P�?      �?                                      �?                                                                              �?      @ui��|��?b�S�	�i?      �?                        	��V��?      �?       @      �?                       @       @               @              �?        �:��?*�H���?              �?      �?        Zas �
�?      �?       @      �?                                               @              �?      �?��>|]�?,�dG��?      �?      �?                              �?                                                                                       @���8�)�?��3��h?                                ���V،?              �?                                       @                              �?       @T�����?4n4s?                      �?        �ԓ�ۥ�?      �?       @      �?       @                               @       @       @                9�)1[��?rM�F�Q�?                      �?      �?!�
���?      �?       @      �?                               @                              �?       @�F���?���{�C�?                      �?      �?      �?      �?       @      �?               @       @       @       @       @       @      �?        m�\d���?b�ދ�g�?                                �@�6�?      �?                       @                                                      �?       @5w\I`��?2md��y�?      �?                        ���Vج?      �?       @      �?               @       @               @       @                      @�����U�?�EQ���?      �?                        ���V،?      �?              �?                                                              �?       @ї�V�i�?����6�?      �?              �?      �?              �?               @      �?      �?      �?      �?      �?      �?      �?              @�U�����?qpTV�?                      �?      �?�@�6�?      �?       @                                                                      �?      �?��<݌�?g�&
�?                      �?        Zas �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �k�.M��?�)��R��?                      �?      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @n��W�?X+���?      �?              �?      �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?              �?       @1[�yj�?`����i�?                      �?      �?�z2~���?              �?               @                       @                       @              @�������?�y�{y�?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�d�Q�ϐ?�9�(� ?                              �?{2~�ԓ�?      �?                       @                       @       @                      �?      �?ٙ�ǰ2�?T^1��?              �?                >�]���?      �?       @      �?       @       @       @               @       @      �?               @=P9��_�?�Z3F��?      �?      �?                              �?       @      �?                                                              �?       @�ئ�N�?��e`��z?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @#w\I`ޓ?�z2P]ǈ?      �?              �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�፿Po�?���Rb�?      �?      �?                �]�����?      �?       @      �?                                       @                      �?       @<��u�4�?���u���?      �?                        3~�ԓ��?      �?       @      �?               @                               @      �?              �?��ǰ2��?�f��q�?      �?                        ��.�d��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�U�����?��k���?                      �?        6���?      �?       @                       @               @                       @      �?      �?Ήo���?偯9��?                      �?      �?[as �
�?      �?       @      �?                       @       @       @       @              �?       @3��x�]�?GB����?              �?      �?        ���.�d�?      �?              �?       @       @       @                       @      �?                rv��?�R�fa��?                      �?      �?�'�K=�?      �?       @                       @                                                       @HT�n��?��2pI�?      �?                        p�z2~��?      �?                                               @                              �?      �?��x�]��?ߝoڊy�?      �?              �?      �?P�o�z2�?              �?               @       @                       @              �?              @q%�yO��?���]��?      �?                        ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                        ����'t�?U��T��?                                ?���@��?      �?       @      �?       @                                                      �?       @��̱���?:��{Vɡ?      �?              �?      �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?               @�d�Q�ϐ?�{Ԃ��?                                ���@��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�፿Po�?���_��?      �?                      �?$Zas �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @)g��1�?-���&�?      �?                        �]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�'�F7�?��:}�?                                P�o�z2�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �6��w�?g[���?              �?                ��Vؼ?      �?              �?                       @                                              �?���I�:�?���-F�?              �?      �?      �?3~�ԓ��?      �?       @      �?                       @               @                      �?      @Q��'�F�?E퐷�@�?                                              �?              �?                                                                      @�/�����?�t�Y=�x?              �?                �D+l$�?      �?       @      �?               @       @               @       @              �?       @�����U�?Nfn�:��?      �?              �?      �?p�z2~��?      �?       @               @       @       @       @       @       @       @      �?      @]�F�?���Z���?                                v�'�K�?      �?       @               @       @       @       @       @       @       @      �?      �?�^!ї��?��"����?      �?      �?                $Zas �?      �?       @      �?                                       @       @              �?        �:��??*i�W��?      �?      �?      �?              �?      �?       @      �?       @       @       @       @       @       @              �?      �?�T�&#�?>���ʲ�?                                �@�6�?      �?       @      �?               @       @       @       @       @              �?      �?Ͽk�.�?uhc~8�?                                              �?                                                                              �?      @�����9�?���W�i?      �?                        ���V؜?      �?              �?                       @       @       @                      �?      @�p��R�?A:	>��?                      �?      �?�@�6�?      �?                       @       @                                                      �?������?��̈́y�?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�d�Q�ϐ?�9�(� ?      �?                        H���@��?      �?              �?                                                                      @Y�ڙ���?�B���?      �?              �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @                ���@��?oؓ [�?      �?              �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�'�F7�?���yӷ�?                      �?      �?�'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @��N�Ա?\Gɶ�7�?      �?      �?      �?        ��V��?      �?       @      �?       @                               @       @      �?      �?       @��¯�D�?�|�V̓�?                      �?      �?P�o�z2�?      �?       @      �?       @               @       @       @       @       @      �?        $X~PT��?��6��?              �?                H���@��?      �?       @      �?       @       @                       @       @              �?      @�V�i���?Q�qhف�?      �?              �?      �?      �?      �?       @               @       @       @       @       @       @       @      �?        d�Q���?֎�����?      �?                      �?              �?                                               @               @              �?      @!s�g�L�?��O��Bs?      �?      �?                ��Vؼ?      �?                                               @                                      @��̱���?]�ZZ�?      �?                        ���V؜?              �?               @       @                                              �?      @���C��?6�
e�΄?              �?                ���V،?      �?              �?                                                              �?        ��6���?�*�ل��?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?8�]�FR�?��ͧ'd�?                      �?      �?���V؜?      �?              �?                                       @                      �?       @�AQ�s��?���M��?              �?      �?      �?v�'�K�?      �?       @      �?               @       @               @       @      �?      �?       @ߚ ���?�fVp�`�?      �?      �?      �?        6���?              �?                       @       @                       @              �?       @�����9�?�1s�p�?                                ���Vج?      �?                       @                       @                                       @�
����?�8���?                                �z2~���?      �?       @      �?       @                                                      �?       @L���S�?�ȅ�ֺ?                                              �?              �?                       @               @       @                       @�FR,?�?7�3��݁?      �?              �?      �?�
��V�?      �?                       @       @               @                       @                (-���?W"�l \�?                      �?      �?�z2~���?      �?       @               @       @       @       @       @                              @���[�?z�%�H�?                      �?        �@�6�?      �?       @      �?       @               @               @       @              �?       @�� Q�E�?z�/HC��?      �?              �?        (�K=�?      �?       @               @       @       @       @       @              �?                )�tN|x�?ۅ�{�X�?      �?              �?        ,l$Za�?      �?       @      �?       @               @                                      �?      �?y4��0�?q�i�u��?      �?              �?        �]�����?      �?              �?                       @               @                      �?        �����?����?      �?              �?      �?�K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @                t+�oM�?�0j.��?      �?                      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����[�?-�CZ���?                                ���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?                F��1��?*�r��?                                              �?               @      �?      �?      �?      �?      �?      �?                      �?�%��}�?����?              �?      �?              �?      �?       @               @       @       @               @       @       @      �?      �?�W���?��ј���?                              �?H���@��?              �?               @                       @                       @                ^�(Ţe�?nm�'�c�?      �?              �?        �ԓ�ۥ�?      �?                       @       @       @       @       @       @       @      �?      @��a�(�?������?      �?              �?        Zas �
�?      �?       @               @               @       @               @       @              �?k� 6\.�?e�� �d�?      �?              �?        ��V��?      �?       @      �?       @               @               @       @              �?       @�N��b�?�i����?                      �?        �RO�o��?      �?              �?       @                       @       @       @       @      �?       @��.h#�?�� ���?                      �?              �?      �?               @      �?      �?      �?      �?      �?      �?       @                �፿Po�?�y!�O��?                                P�o�z2�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?���@��?�i�����?      �?                        ���V،?      �?              �?               @                                                       @S,ZV��?��y�ek�?                      �?      �?�z2~���?              �?               @                       @                      �?              �?��+$��?�:�n*�?      �?              �?      �?e�v�'��?      �?       @                               @                       @       @              �?��l��?�:��	�?              �?                �'�K=�?      �?                       @               @       @       @               @                �bѲ
n�?4��h�l�?                                �V�H�?      �?              �?                       @                                      �?      �?	�{B��?�np���?      �?      �?      �?        �'�K=�?      �?       @                                                                      �?       @���-�<�?��5vl�?      �?                        6��9�?      �?                                                                              �?        �{'Y��?
4)��?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @                F��1��?���F�	�?      �?                      �?��RO�o�?      �?              �?       @       @       @                       @      �?               @q��3���?.�n����?      �?              �?              �?      �?                       @       @               @       @       @       @      �?        d��ht�?�g��,�?      �?              �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @                �U�����?A:	>��?                                �
��V�?      �?                               @       @                       @       @      �?      @�1����?��W����?                      �?      �?H���@��?      �?                               @       @               @       @      �?              �?�|�?^�?�	��?                              �?���V؜?      �?                       @                       @               @              �?        F��s�?j�寚��?                                �RO�o��?              �?                       @                       @       @              �?       @]<��u��?M�Y�8�?                              �?�z2~���?      �?                                                                              �?       @�9�፿�?�A0��H�?      �?                                      �?                                                                              �?      @���"X~�?U�9��g?      �?              �?      �?	��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @qi��|��?4��+D�?                                ���V،?              �?                                                       @              �?       @Sb����?�8S]f�t?      �?              �?      �?P�o�z2�?      �?                                       @       @       @       @       @      �?        �}��j�?~���8�?                      �?        ��V��?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?uhc~8�?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @�����`�?d��]�a?                                              �?                                                                                      @ꏗ�(��?��ׇh?      �?      �?                ���V؜?              �?                               @                       @              �?       @S��*�?�Ms�̊?                                �D+l$�?              �?                                       @               @      �?      �?      �?�S��%�?�}7gA�?                                ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�m��W�?��	���?      �?                      �?��.�d��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?Rp�l?�Bt�n�?      �?                        ��V��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        \��r�?�qhف3�?                              �?���V؜?      �?                       @                       @                              �?      @xwwwww�?��^l�?      �?                        �K=��?      �?                       @               @                              �?              @�:��?��T���?                      �?        ���.�d�?      �?       @      �?       @               @               @               @      �?      �?�q%�yO�?x�S���?      �?                      �?              �?               @      �?      �?      �?      �?      �?      �?                      @nC��x�?��q�S~-?      �?              �?        Zas �
�?      �?       @               @               @                       @       @      �?      @X-�r�?6�k-|�?      �?                                      �?       @                               @       @                                      @Z�KS}��?�?93qt?              �?                ���V،?      �?              �?                                                              �?       @�l	�Y�?�7�!\��?                                 �
���?      �?       @      �?                                                              �?        S,ZV��?��*o@��?                                �'�K=�?      �?       @      �?                                       @       @                        �:��?я��&n�?                                �D+l$�?      �?       @       @      �?      �?      �?      �?      �?      �?       @               @h#���?�g?ʤ��?                      �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @              �?�2��?.�H���?                                �'�K=�?      �?                               @       @       @       @               @              @����e�?����<��?      �?                         �
���?      �?       @      �?                               @                              �?       @�~5&��?w����?                                ���V،?      �?              �?                       @                       @              �?      @�a�(Ţ�?������?                      �?      �?�ԓ�ۥ�?      �?              �?       @               @       @       @       @              �?       @]I`�:�?�AYm��?      �?              �?      �?��RO�o�?      �?                               @               @       @                              �?I!�i��?W&s���?      �?      �?      �?        F���@��?      �?       @      �?       @       @                               @              �?      �?c9�W�?�Y=�T�?              �?      �?        ,l$Za�?      �?              �?       @       @               @                              �?       @Ͽk�.M�?������?      �?                        ��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              @E�(Ţe�?<q��ҳ?                                >�]���?      �?       @      �?       @       @                       @       @              �?      �?Ɉ���!�?A֬�̱�?                      �?        ܥ���.�?      �?              �?               @       @               @       @      �?      �?       @5A .�?�Z>�}B�?              �?      �?        3~�ԓ��?      �?       @      �?               @       @               @       @              �?       @�mZq�$�?��.J:��?      �?              �?      �?      �?      �?       @      �?       @       @       @       @       @       @       @                �w�ӥ��?$d�_���?              �?                v�'�K�?      �?       @      �?               @                                              �?      �?*L����?̫�8�?      �?      �?      �?      �?�V�H�?      �?       @      �?       @       @       @               @                      �?       @��S�@�?�R�\
��?      �?                        Zas �
�?      �?                                               @                              �?      @5w\I`��?�3��4�?      �?              �?        ��ۥ���?      �?       @      �?       @       @       @               @       @      �?      �?       @�D)�?y������?      �?              �?        ��ۥ���?      �?       @      �?                                       @       @              �?       @r@���?x��̈́�?                      �?      �?      �?      �?       @               @       @       @       @       @               @                ZV����?��ߧ��?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      �?���@��?�v)k���?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?                        ��N�ԑ?�]Q�T�?              �?                 �
���?      �?       @      �?               @                       @                      �?       @��Y;��?��F����?                      �?      �?�z2~���?      �?                       @               @       @       @       @       @      �?      @�����?�V���?      �?                      �?�'�K=�?      �?       @               @       @       @       @       @       @       @              @�r�9ֳ�?�]V�kp�?      �?              �?      �?��ۥ���?      �?       @      �?               @       @               @       @       @      �?        �*g���?�ɡxs�?                                ���Vج?      �?                       @               @                                              �?ͤ=����?�9�(��?      �?                        �V�H�?              �?               @               @       @       @       @       @      �?        �w����?W1�!�:�?      �?                        �'�K=�?      �?       @      �?                                                              �?      @T�n�Wc�?�V"�l�?                      �?      �?���.�d�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @���Z��?�d��?      �?              �?        �'�K=�?      �?              �?                                                              �?        ���&�?��V��?      �?                        �V�H�?      �?       @      �?       @                               @                      �?      �?��Y;��?�Q�}7�?                                ���Vج?      �?                                                                              �?      �?�bѲ
n�?����H��?      �?              �?      �?�ԓ�ۥ�?      �?       @                                       @       @       @      �?      �?        ui��|��?�� ���?                                              �?       @      �?                                       @                      �?       @l	�Y �?w�\�?                                �V�H�?      �?       @      �?       @       @                                                      @~5&��?�>���F�?                      �?        �z2~���?      �?                       @                       @                                        �
����?s�e̮׳?      �?                        �
��V�?      �?       @      �?               @       @               @       @              �?       @Gm?C��?U�Y"���?                                              �?                                                                              �?      @�r@��?EF�=?h?                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?^��Z��??ښo;�?                      �?      �?�o�z2~�?      �?              �?               @       @               @       @              �?       @w\I`��?:i׊�!�?      �?                        ��Vؼ?      �?       @      �?                                       @                      �?       @%K!�i�?�QF! ն?              �?                              �?              �?                                       @                               @��I{+�?�iiǔ1|?                      �?      �?$Zas �?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      @)���O�?#�Blv�?                                [as �
�?      �?                               @       @       @       @       @       @              @��.h�?�)�M�?                      �?      �?��RO�o�?      �?              �?                                                                       @��6���?�9�[�?                                {2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        M:'>��?XT�9�?      �?                        ���V،?      �?              �?                       @                       @              �?       @z�Τ=��?��r��?                                ��V��?      �?                       @       @               @                       @      �?      @��U�?<(��z�?                                �K=��?      �?       @      �?       @       @       @               @       @              �?      @�9ֳv&�?)�6T�Z�?                                �'�K=�?      �?       @               @       @               @                                      @�����T�?�.]�AS�?      �?              �?        6��9�?      �?       @      �?                       @       @       @               @              @J�hY7�?�'A��k�?                      �?      �?{2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?       @                ����[�?���zh�?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?����[�?ό2
��?      �?              �?        Zas �
�?              �?               @               @       @       @       @       @      �?      @e�����?�6����?      �?      �?              �?�6��?      �?       @      �?       @                                                      �?      @*L����?0؈��7�?      �?                        �K=��?      �?       @      �?               @       @               @       @              �?       @����>�?����?      �?                        F���@��?      �?              �?                                               @              �?       @B�/����?�Ҟ>�?                      �?      �?6���?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?Xph>ׯ?{�M%���?                      �?        ��ۥ���?      �?       @                               @       @       @       @       @      �?        *L����?L�*����?      �?                        ���V؜?      �?              �?       @                                       @              �?      @�����?.�{��?              �?                ���V،?      �?       @                       @                                              �?      �?�g�L�c�?��.骀�?      �?              �?      �?e�v�'��?      �?              �?               @               @                       @      �?        �`�AQ��?ɳ�y�	�?      �?                        6��9�?      �?              �?       @       @       @               @       @              �?       @A���Kn�?�)��6d�?              �?      �?              �?      �?       @      �?               @       @       @       @       @       @      �?      �?����w�?��X	�?              �?                              �?              �?                                                              �?       @�7�B�]�?���x?      �?              �?      �?(�K=�?      �?       @               @       @       @       @               @      �?                &`��"�?�0\�M
�?      �?      �?              �?�@�6�?      �?                               @               @                              �?       @�
n���?�k=r�4�?                                              �?              �?                                       @                               @�G��q
�?U�B.|?      �?              �?      �??���@��?      �?       @      �?                       @               @       @                       @�3i�ae�?���U��?                                ?���@��?      �?                               @                                                      �?Q,?(��?B;�m,P�?                                              �?                                                                              �?      �?�9�፿�?��Y�pWh?      �?                      �??���@��?      �?                       @                                                               @*L����?������?                      �?        �ԓ�ۥ�?      �?                       @                               @              �?      �?        e�����?�O�u 9�?      �?                                      �?                                                                                      @�?���}p�h?                      �?        ���V؜?      �?       @      �?                                                              �?      �?]�;x��?�t�Y=��?      �?      �?      �?        6��9�?              �?                       @       @                                      �?      �?���7q�?��J{~�?      �?                        ��V��?      �?              �?               @       @                                      �?      �?T�n�W�?!ad1,��?                              �?���Vج?      �?                                               @                              �?      @w�����?�^,5쪟?      �?              �?        �ԓ�ۥ�?      �?       @      �?                                                              �?       @��g{�?\�TQ��?      �?              �?        ��V��?      �?       @      �?               @                       @                      �?        �፿Po�?_�n"��?      �?              �?      �?SO�o�z�?      �?       @      �?       @                               @       @      �?               @��vA�?[u�X���?      �?                        �]�����?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �'�F7�?��?�?                      �?      �?H���@��?      �?       @      �?                                       @       @              �?        r@���?������?      �?      �?                P�o�z2�?      �?       @      �?               @       @                       @              �?       @�	�p��?9��չ��?              �?      �?        ��.�d��?      �?       @      �?       @       @       @               @       @              �?       @�"s�g��?j�OA��?              �?      �?        �RO�o��?      �?       @      �?               @       @               @       @              �?       @r@����?.�+Z��?      �?              �?      �?      �?      �?       @      �?       @               @               @       @       @      �?        ��+	��?�po����?      �?              �?      �?P�o�z2�?      �?              �?       @               @                               @              �?���!���?��V`��?                      �?        �K=��?      �?       @      �?               @       @               @       @      �?      �?        Gm?C��?kZ�P�?                      �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ����[�?�P-�2�?                              �?	��V��?      �?       @                               @                              �?      �?      @V:'>���?��<�#�?      �?      �?                ���V،?      �?                       @               @               @                                �w�ӥ��?�����?      �?                        �z2~���?      �?       @      �?       @               @       @       @       @              �?      �?��l��?��b`C�?              �?      �?        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�X����?o.����?      �?      �?      �?        (�K=�?      �?       @      �?               @       @               @       @      �?      �?       @Y7���?� �yg��?      �?              �?      �?[as �
�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�rv��?YMM2�õ?      �?      �?                ���V؜?      �?       @      �?               @       @               @       @              �?       @e0
84��?X)�*I�?                                ���V؜?      �?       @      �?                                                              �?       @���I�:�?���Kdؗ?                                �@�6�?      �?       @      �?       @                                                      �?        T�n�W�?���0��?                      �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @\��r�?A]��3�?                      �?      �?H���@��?              �?               @       @       @               @       @              �?      �?,ZV���?����?                      �?              �?      �?       @      �?       @       @                               @       @      �?      �?�Gm?C�?�!w�U}�?      �?                        ��RO�o�?      �?              �?                       @                                               @0�	��?�^ۛ:�?      �?              �?      �?H���@��?      �?       @       @      �?      �?      �?      �?      �?      �?              �?        ���6�?a���2�?              �?      �?        �@�6�?      �?              �?                               @       @                      �?       @�dsǕ�?1pI$q�?      �?                                      �?       @               @       @                                                       @�#�d�Q�?�j�Mt?              �?      �?        P�o�z2�?      �?       @      �?       @       @                               @      �?      �?      �?�Up�l��?�ʟ<�?                      �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @                �d�Q�ϐ?��o�W>�?      �?              �?        ��RO�o�?      �?       @      �?       @               @                       @                       @1[�yj�?��<Y��?      �?              �?        ��RO�o�?      �?       @      �?               @       @                                      �?       @�%��f��?T�զ9�?                      �?        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                      @9�%��}�?��{#%y?                      �?        �@�6�?      �?              �?               @       @       @                      �?      �?        �a�(Ţ�?���I��?      �?              �?        �D+l$�?      �?       @               @                       @               @      �?      �?      @%�yO�0�?%ꘓ�?                      �?              �?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?)g��1�?��}M"	�?      �?                        v�'�K�?      �?       @       @      �?      �?      �?      �?      �?      �?      �?                n��W�?���I���?              �?      �?        SO�o�z�?      �?              �?       @                                                      �?      �?!�����?|)�����?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�X����? �<$3?                      �?        Zas �
�?              �?                                       @       @       @              �?       @uN|x�/�??����`�?                      �?        �z2~���?      �?              �?                               @       @       @       @      �?      �?��a��?B��M8��?                              �?H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?����'t�?jQV��?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?       @              @��N�ԑ?#"�b�a�?                      �?        ��ۥ���?      �?       @               @       @       @       @       @       @       @              �?�@��~�?A������?      �?              �?        SO�o�z�?      �?       @               @                       @       @       @      �?              �?*L����?�U�����?              �?      �?         �
���?      �?       @      �?               @       @                       @              �?       @m��W�?��s�?                                      �?      �?       @      �?       @       @       @       @       @       @       @      �?       @P_W-��?Y��;0N�?      �?              �?      �?���Vج?      �?               @      �?      �?      �?      �?      �?      �?      �?               @�፿Po�?
��IG�?                      �?      �?�@�6�?      �?       @      �?       @       @                       @                      �?        J�hY7�?�`�P���?      �?      �?      �?        ��ۥ���?      �?       @      �?                                               @              �?      �?UUUUUU�?��CmA��?      �?                                      �?              �?                                                              �?       @���U�?�^��w?                                F���@��?      �?       @      �?       @                               @       @              �?       @���+$�?����?                                �z2~���?      �?       @      �?                       @       @                              �?       @���[��?��/~���?      �?                      �?              �?              �?                                                              �?       @�=�� �?m[����x?      �?                        �]�����?      �?       @      �?               @                                              �?       @d��ht�?l����G�?      �?                        �@�6�?      �?                       @               @       @       @       @       @      �?      @!�iŽ�?,'ʬA
�?      �?                        �@�6�?      �?              �?               @               @       @              �?      �?       @�r�9ֳ�?g!ի�g�?                      �?      �?���V؜?      �?              �?               @               @                              �?       @M+�d��?Ef��J�?                      �?        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�]�FR�?��,�p��?                      �?      �?!�
���?      �?       @      �?                       @                       @      �?      �?       @�
����?������?                                              �?                                                                                      @6��`�A�?f��	i?                      �?      �?�@�6�?      �?                       @       @               @       @       @       @               @��I{+�?�p�AX��?      �?                        �V�H�?              �?                       @                                                        ��̱�?�K�]�?              �?      �?                      �?              �?                                                              �?      @��J��?d�g$�ix?      �?      �?                �ԓ�ۥ�?      �?       @      �?       @                                       @                      �?�jL�*�?ƫ�4�Y�?                      �?        H���@��?      �?                       @       @               @               @              �?      @�d�Q���?�1�h���?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?              �?       @�d�Q�ϐ?�9�(� ?                      �?      �?���V؜?      �?       @                       @       @               @                      �?        �Kn��4�?u�N����?              �?      �?      �?Zas �
�?      �?       @                               @               @              �?      �?       @dsǕ��?`����$�?                                ?���@��?      �?               @      �?      �?      �?      �?      �?      �?                      �?1[�yj�?���E~?      �?      �?      �?        �D+l$�?              �?               @               @       @       @       @       @      �?      �?S��*�?�;�X���?      �?                        ���V،?      �?              �?                       @               @       @              �?       @�>|]��?��Mc�#�?                                 �
���?      �?              �?       @               @       @                      �?      �?      �?Ln��4��?�tE���?      �?              �?        �D+l$�?      �?       @      �?                                       @       @              �?      �?z����"�?���t��?                      �?      �?              �?              �?                                                              �?       @ї�V�i�?:j)��x?      �?                        ?���@��?      �?              �?                                               @              �?       @ȕ�=��?����?      �?              �?      �?      �?      �?       @               @       @       @                               @              �?��Ͽk�?\�܌\�?      �?              �?        ���V؜?      �?       @      �?                               @                              �?        ��<݌�?d������?                      �?        ��RO�o�?      �?       @               @                               @                      �?        &��f���?o�g,>�?      �?                      �?�@�6�?      �?       @      �?       @                                                               @���!���?,�>s��?      �?              �?      �?�ԓ�ۥ�?      �?                       @               @       @       @       @                       @ئ�N��?�<���?      �?              �?      �?Zas �
�?      �?                       @       @       @       @       @       @      �?                 ʣ��8�?l�)K�^�?                      �?        �D+l$�?      �?       @      �?               @                       @       @                       @�ht3Na�?���M�;�?      �?              �?        �D+l$�?      �?       @      �?                       @               @       @      �?      �?        �۴���?�K��F��?                      �?      �?�'�K=�?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @O�)���?IF��/�?      �?                        ��RO�o�?      �?                       @                                                              @���7q�??�q����?      �?              �?        �RO�o��?      �?       @      �?               @       @               @       @      �?                I�:Bl��?i��n��?      �?      �?                $Zas �?      �?              �?                                       @       @                       @��7q��?@Z�'�?      �?              �?        ,l$Za�?              �?                       @       @               @       @       @                ����?Q0�ۃ�?                                �6��?      �?       @               @       @       @                                      �?        [�<��?Z��R}�?      �?      �?                �@�6�?      �?              �?                                               @              �?       @ph>�/�?PEV��D�?      �?              �?      �?���Vج?      �?       @      �?       @               @                                      �?       @�s��2�?p�V���?      �?      �?                ��Vؼ?      �?       @               @                                                               @�
n���?��qs�?      �?      �?      �?      �?��V��?      �?       @      �?       @       @                                              �?       @�@��~�?_j7���?                                [as �
�?      �?       @      �?                                                              �?       @�c=kg�?b���YP�?      �?                        ���Vج?      �?              �?                                       @                      �?      @���U���?��5��o�?                              �?              �?                       @                       @                                       @,u�ئ�?~�i���p?                                ���V؜?      �?       @                                       @       @                      �?       @��-��?h�K�+�?                      �?              �?      �?       @      �?       @       @       @       @       @       @       @      �?        t�ئ��?m6�L��?      �?                         �
���?      �?                                               @       @              �?              �?H���<�?�/��3��?      �?      �?      �?        {2~�ԓ�?      �?       @      �?       @                               @       @                       @aJ̖p��?���9
�?      �?                        F���@��?      �?              �?       @                                                              @,�����?{-�Fj�?      �?                      �?	��V��?      �?                                                                      �?              @X�ڙ���?�>�]ݒ�?                                $Zas �?      �?       @                       @               @               @              �?      �?V�ߚ �?�rV���?      �?              �?      �?�RO�o��?      �?       @      �?       @               @               @              �?      �?        r@���?�A�Ud�?                      �?      �?Zas �
�?              �?                       @       @       @       @       @       @      �?        �X����?�J%,h��?      �?              �?        �RO�o��?      �?                       @                               @              �?      �?      @�^<��u�?~��1)�?                                [as �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�L�5A �?�	ok�γ?                      �?        6���?              �?               @       @                       @              �?      �?       @6��`�A�?99��ɞ�?      �?                                      �?              �?                                       @                      �?       @�?^���?�g�D��|?      �?                      �?v�'�K�?      �?                               @       @       @       @       @       @      �?      �?�?^���?^qƦ�?                      �?      �? �
���?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�U�����?	0��� �?                      �?      �?���.�d�?      �?       @      �?               @       @       @       @       @      �?      �?       @�\d����??�|����?      �?              �?        3~�ԓ��?      �?                       @       @               @       @              �?              �?o��z��?��Ʊ[�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?              �?      @nC��x�?@Ր�,?                      �?      �?�ԓ�ۥ�?      �?       @      �?               @       @       @       @       @      �?      �?        ���(���?�w@o��?      �?                        [as �
�?      �?       @      �?               @                                              �?       @*L����?@g���?              �?                v�'�K�?      �?       @      �?       @                               @       @       @      �?        � Q�E��?s5��?              �?      �?        SO�o�z�?      �?       @      �?                                       @       @              �?       @����'t�? �����?                                              �?                                                                                       @�vAIE�?�:�:�g?                      �?        �'�K=�?      �?               @      �?      �?      �?      �?      �?      �?                        ����[�?�$)��=�?      �?                        	��V��?      �?       @      �?       @       @       @       @       @                      �?        �S��%�?ap9#{k�?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @                �U�����?�D�}�U�?      �?      �?      �?        3~�ԓ��?      �?       @      �?                                               @              �?       @�_���@�?QqJ�_�?      �?                        6���?      �?                               @       @       @       @               @                cX�~k��?��t�m��?      �?                        �z2~���?      �?       @      �?                       @                                      �?       @�����?@�9��	�?      �?              �?        ��ۥ���?      �?              �?       @                               @       @              �?       @��R���?�ʌU��?              �?                �z2~���?      �?       @      �?                       @                                      �?      @d��ht�?�#;���?      �?              �?      �?�'�K=�?      �?              �?                                                              �?       @L�*g��?Iw���?      �?              �?      �?!�
���?      �?       @      �?               @               @                      �?                T�@ʾ��?\�M
���?                      �?      �?�z2~���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?��N�Ա?Ki���<�?                              �?,l$Za�?      �?       @                       @                       @       @      �?      �?      @�[���?�h�C�~�?      �?                        6��9�?              �?                                               @               @              �?�R,Z�?%��d,�?                                ���V،?      �?       @      �?               @                                                       @q
Sb���?��y�ek�?                                �]�����?      �?                       @                                                      �?       @፿Po�?nc��0o�?                              �?�V�H�?      �?       @      �?                       @       @                              �?        y4��0�?�p��?      �?                        �z2~���?      �?       @      �?                                                              �?       @S,ZV��?յd�}��?      �?                        $Zas �?      �?       @               @                       @                                        x\I`��?���`Q�?      �?                        P�o�z2�?      �?              �?               @       @                              �?              �?4�G�Ɉ�?��3���?                                ��Vؼ?      �?                                                                              �?       @o�Wc"=�?��k��ۦ?                      �?      �?��RO�o�?      �?              �?               @               @               @              �?      �?h{����?i�/k��?                      �?        (�K=�?      �?       @      �?                       @       @       @       @       @      �?        ��0%f�?�oڊy�?      �?              �?      �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�%��}�?kz'��?                      �?        �'�K=�?      �?       @                                                                      �?       @��x�]��?�2��s�?                                ��V��?      �?              �?                                                              �?        �V�ߚ�?B�K.r��?      �?      �?      �?        �'�K=�?      �?       @                       @       @               @              �?      �?      �?�/�����?��Y-�o�?      �?                        SO�o�z�?      �?       @      �?                       @                                               @ȕ�=��?�gg1�T�?                      �?      �?���Vج?      �?                                                                                      @q%�yO��?G�0��ӗ?                                �ԓ�ۥ�?      �?       @      �?       @       @       @       @       @       @       @      �?      @e� �;�?�Bc��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                        F��1��?��ֺ�?                      �?      �?ܥ���.�?      �?       @      �?                                               @      �?      �?      @��"X~P�?�K����?                                              �?               @      �?      �?      �?      �?      �?      �?                      @���@��?�ppTV�)?                                ���Vج?      �?                       @                       @                                      �?[ݧ����?��3.z�?              �?      �?        �RO�o��?      �?       @      �?                       @               @       @      �?      �?      �?����e0�?�Q|�v1�?                                3~�ԓ��?      �?       @      �?       @               @       @       @       @      �?      �?        �C��?}'�;ā�?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              @F��1��?�t���`�?      �?              �?      �?�'�K=�?      �?                       @                                       @              �?      @�
����?"��
:��?      �?                        ��ۥ���?      �?       @      �?                                               @              �?       @ ʣ��8�?�d��S��?      �?                        6��9�?      �?       @      �?                                               @              �?        �6��w��?�:o[�?                      �?      �?p�z2~��?      �?       @               @       @       @                               @               @w�D_r[�?5o�����?      �?                        �6��?      �?       @               @       @       @       @                                       @��j1v�?ļ���|�?                      �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                \��r�?��?l�)�?                      �?        �
��V�?      �?       @      �?               @       @               @       @              �?      �?��8�)1�?i�u�b��?                      �?        �ԓ�ۥ�?      �?              �?                                                              �?       @p�l�?Ȋ��3��?                      �?        {2~�ԓ�?      �?       @      �?       @               @               @       @      �?                �b�V��?�Ģ���?      �?                                      �?              �?                                                              �?       @p�l�?��Y�pWx?                      �?        ܥ���.�?              �?                       @       @                              �?              @Sb����?�?.��k�?      �?              �?        �@�6�?      �?                                                       @                      �?        �፿Po�?����h�?      �?              �?      �?��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �X����?�ع�(7�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @m+�oM�?V�I�?              �?      �?              �?      �?       @      �?       @                                               @                ph>�/�?$����?                      �?        �@�6�?      �?       @      �?       @       @       @       @       @       @              �?        |k� 6\�?��$����?      �?                        �ԓ�ۥ�?      �?       @               @       @       @       @       @       @       @              @�ߚ ��?'���F�?      �?                        ?���@��?      �?                                                               @              �?      @��W��?��"����?                      �?      �?��RO�o�?      �?       @      �?                       @                       @              �?       @���[��?��n��O�?      �?              �?      �?6��9�?      �?              �?                                       @       @      �?              �?	�U:�?~p�L��?      �?      �?      �?        ��ۥ���?              �?               @       @       @       @                       @              �?�@ʾ���?�#k��?      �?              �?      �?F���@��?      �?                               @       @       @                                        �������?=LLg��?                      �?        !�
���?      �?              �?       @       @       @               @              �?      �?       @����?�2����?      �?                      �?�
��V�?      �?              �?       @                                                      �?        �ae��	�?���F�?      �?                      �?���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @���C�?��$�f?                                              �?       @       @      �?      �?      �?      �?      �?      �?              �?       @��+$��?7c��"J?                      �?      �?e�v�'��?      �?                       @               @       @               @       @                ��j1v�?��Rj�t�?      �?      �?      �?        �'�K=�?              �?                                               @       @              �?       @��j1v��?ᗊ����?                      �?      �?�@�6�?      �?                                                                              �?       @�=�� �?�+r�κ?      �?              �?      �?6��9�?              �?               @       @       @                                                h�����?*@��"�?      �?              �?      �?�
��V�?              �?               @               @       @       @              �?              @]<��u��?��_�4�?      �?                        	��V��?              �?                                                                      �?      @g�)L�ٲ?u�J=��?                                �@�6�?              �?               @                       @                       @              @l��4�u�?�E&��3�?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @^��Z��?��?Q��?      �?                        6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�0[�yjv?}�u^Ş?      �?                        �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�]�FR�?�\5ܴv�?      �?              �?      �?�K=��?      �?       @      �?               @                       @       @              �?        �n�)L�?C��%m�?      �?              �?      �?��Vؼ?      �?              �?                       @       @       @       @                       @o��T�?��h���?              �?      �?         �
���?      �?                                       @                       @      �?              @2��g�?s�(:Q�?      �?                        6��9�?      �?       @      �?       @                               @       @                       @��r��?����<�?              �?      �?              �?      �?       @               @       @       @       @       @       @       @      �?        t3NaJ��?��ЯA��?              �?      �?        �K=��?      �?       @      �?       @               @               @       @      �?      �?      �?��>�MF�?���N�?      �?      �?                F���@��?              �?                       @               @               @              �?       @?y4���?�f3­/�?                      �?      �?      �?              �?               @       @       @       @       @       @       @      �?      �?dsǕ��?�/M���?      �?                      �?ܥ���.�?      �?       @               @       @       @                              �?      �?         .�c�?���FG�?                                p�z2~��?      �?       @               @               @       @                       @      �?      @I!�i��?`�17!�?                                              �?               @      �?      �?      �?      �?      �?      �?                      @�m��W�? Ր�,?                      �?      �?�]�����?      �?              �?                                               @              �?       @��̱���?��uq�+�?      �?                        �D+l$�?      �?               @      �?      �?      �?      �?      �?      �?       @              @,1[�yj�?�Ea�x�?      �?                        ��Vؼ?      �?       @                                                       @                      @Ήo���?�H��_�?      �?              �?        3~�ԓ��?      �?       @                               @       @       @       @       @              �?A .��?�����?                                ���V،?      �?                               @                                              �?      @�7q���?r	婆?      �?                        ��RO�o�?      �?                                       @                       @      �?      �?       @d����I�?cH����?      �?                        ���V،?      �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?'�d��+\?      �?              �?      �?�ԓ�ۥ�?      �?       @      �?               @       @       @       @       @              �?       @ۙ�ǰ2�?�A8}��?                      �?              �?      �?       @      �?       @       @       @               @       @       @      �?      �?��Ͽk�?�� !���?              �?                              �?              �?                       @                                      �?        ���H*�?sn:Oo�z?                                �z2~���?      �?              �?                       @       @               @              �?       @��%���?��ٷ�Ͽ?      �?              �?      �?6���?      �?       @      �?               @               @       @              �?      �?      �?c9�W�?�w`����?                      �?      �?��ۥ���?      �?              �?                       @                               @               @�c=kg�?Q��R�?      �?                        ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?���'th?�|�V̳?                      �?        {2~�ԓ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�]�FR�?����F}�?      �?      �?      �?        ��V��?      �?       @      �?               @       @               @       @              �?       @}䛌8j�?@Fg\�8�?      �?              �?      �?�RO�o��?      �?              �?               @       @               @              �?               @9�WH�%�?��[�X�?                      �?              �?      �?       @      �?       @               @       @       @       @       @      �?      �?�ć7�B�?$��Z�?              �?      �?      �?�@�6�?      �?       @      �?                       @                                      �?      �?V����?�-1��?      �?              �?        6���?      �?               @      �?      �?      �?      �?      �?      �?       @              @nC��x�?/�l>=�?                                �z2~���?      �?       @                                       @       @       @      �?      �?      @
n��W�?�������?      �?                        ���Vج?      �?                       @                       @                              �?      @HT�n��?�FwR�?                                      �?      �?       @      �?                       @       @       @       @       @      �?      �?���-�j�?�yӷ[��?                      �?      �?$Zas �?      �?       @               @                               @       @      �?                T�n�Wc�?y�fQ0�?              �?                (�K=�?      �?       @                       @       @       @       @               @      �?        ���I�:�?ᘶ�-�?      �?                        6��9�?      �?              �?                                                                      @'#��~��?cx���+�?      �?              �?        H���@��?      �?              �?               @                       @                      �?      �? J�hY�?�;�0��?                                ܥ���.�?      �?                       @       @                                       @              �?�#�6���?�Y�(�C�?                      �?      �?P�o�z2�?      �?       @      �?               @               @       @       @       @      �?      �?Wc"=P9�?=�����?                              �?�@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      �?^��Z��?��KS�?      �?      �?      �?        �V�H�?      �?              �?                                               @              �?       @g��}���?8��y|�?                      �?      �?��V��?      �?                       @       @       @                              �?                z�D_r�?h�g�x�?                                �ԓ�ۥ�?              �?                               @       @                              �?       @�����?v�q"}b�?      �?                        �]�����?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?�d�Q�ϰ?,'ʬA
�?                      �?      �?��RO�o�?      �?                       @       @               @                                        H���<�?����?                      �?      �?�o�z2~�?      �?       @      �?       @                               @       @       @      �?        �3i�ae�?�5��{q�?                                �
��V�?      �?              �?               @       @                                      �?       @��'�?��:	��?                              �?v�'�K�?      �?       @      �?       @               @       @                       @      �?      �?9�WH�%�?�������?      �?              �?        ��.�d��?      �?       @                       @               @                                        z�D_r�?�6�t�D�?                      �?      �?3~�ԓ��?      �?       @      �?       @                               @       @      �?      �?      �?�p����?S`(G:<�?                                F���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�d�Q�ϐ?5�? =�?                      �?        SO�o�z�?              �?                       @               @                      �?              @�ti��|�?������?              �?      �?        F���@��?      �?       @      �?                                               @              �?       @�>�MF�?�O4���?                                �z2~���?      �?              �?               @               @                              �?      @��&`�?~�N��?                      �?      �?>�]���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?-h#���?(���~C�?      �?                        �V�H�?              �?               @               @       @                       @              @�C��x�?W�{^D��?      �?              �?      �?Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?       @              @���@��?�E#�-�?      �?                        6��9�?      �?              �?       @       @       @       @       @       @              �?       @$����>�?sҮ�C�?      �?              �?      �?���.�d�?      �?       @      �?       @       @       @                                      �?       @.�c=k�?m������?              �?      �?        �
��V�?      �?       @      �?               @       @       @       @       @              �?       @���>|�?�3����?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                       @����'t�?�G�O��?                      �?      �?�]�����?      �?               @      �?      �?      �?      �?      �?      �?      �?              @��N�ԑ?!4����?                                e�v�'��?      �?       @      �?                               @       @       @              �?       @��T��?\e����?              �?                $Zas �?      �?              �?                                       @                                �AQ�s��?�g�x���?      �?                        ?���@��?      �?       @      �?               @                                                       @��I{+�?�.���c�?      �?              �?      �?��V��?      �?                       @                       @       @       @       @      �?        	�{B��?$�}����?              �?      �?      �?�
��V�?      �?       @               @               @       @       @              �?               @#�6��w�?T����?      �?              �?      �?��.�d��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @I`�:�?=R���a�?                                P�o�z2�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�X����?g�<��?              �?                ?���@��?      �?              �?               @       @               @       @              �?      �?!ї�V��?�b
��?                      �?      �?�]�����?      �?       @      �?                       @               @       @              �?        ��E���?��6A���?      �?      �?                                      �?                               @                       @              �?       @���vA�?��ᦵc?      �?                        6��9�?              �?                                                       @              �?      @@�/����?ABy���?      �?                        ?���@��?              �?                                       @               @              �?       @=Q�s���?�:��^��?                                Zas �
�?      �?       @      �?                                                                       @C�]�FR�??H�%�\�?                                      �?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����`�?f;=����?              �?      �?        e�v�'��?      �?       @      �?       @       @       @       @       @       @      �?      �?        ��^<��?�o�����?      �?      �?                ��V��?      �?              �?               @       @               @       @              �?        u�4�G��?[I���?                      �?      �?���@��?      �?              �?                       @       @       @       @      �?              @�L�5A �?on�����?      �?              �?        �ԓ�ۥ�?              �?                       @       @       @       @       @      �?      �?      �?>|]��?%���X�?              �?                >�]���?      �?       @      �?               @       @       @       @               @      �?        �f��}��?*Խ�i �?                                                      �?                                                                      �?      @qi��|��?G,˽H?      �?              �?      �?(�K=�?      �?                       @       @       @               @       @       @      �?      �?��̱���?*����?                      �?        �D+l$�?      �?       @      �?       @       @                       @                      �?       @&���[�?=/"Ӵ��?      �?              �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @M:'>��?�r���ճ?                      �?        6��9�?      �?       @               @               @       @                      �?              �?�S�@ʾ�?��uq�+�?                      �?      �?�]�����?      �?                               @               @                                       @�a/��?��8
?��?      �?                                      �?              �?                                               @                       @�~5&��?S�.��)}?      �?      �?      �?        �
��V�?      �?       @      �?               @               @       @       @              �?       @��V�i��?�d} �?      �?                        �
��V�?              �?                                       @                              �?      �?��a/�?�p)-�e�?      �?                        ��.�d��?      �?                       @               @                              �?               @N��b��?v��zx�?                                ��RO�o�?      �?              �?               @               @                              �?      �?���w��?$����&�?      �?      �?      �?        Zas �
�?      �?       @      �?                                       @                      �?      �?H*��E�?���!&E�?                      �?      �?$Zas �?      �?                       @                                                              �?�'�F7��?di���<�?                      �?      �?�@�6�?      �?                       @                                                                w�����?<��䠰?                      �?      �?�ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @�rv��?�wx��?      �?              �?      �?6���?              �?               @       @       @               @              �?              @��e0
8�?��;Ͼl�?                                �K=��?      �?                       @       @                               @      �?               @w�D_r[�?�|�8��?      �?              �?        [as �
�?      �?       @                                               @                      �?      �?䛌8j��?2���.��?                                �z2~���?      �?       @      �?               @                               @              �?       @��Y;��?�|T�x��?                                ��V��?      �?       @      �?               @       @               @       @                       @E�Ήo�?.�b���?      �?                        F���@��?      �?              �?                                       @       @              �?       @� 6\.2�?�$��<�?                      �?      �?�z2~���?      �?              �?               @       @       @                                       @:]��#��?�4?;*��?      �?                      �?              �?       @      �?                                                              �?       @,�����?��c|Az?      �?                                              �?                                                       @              �?        �,u�ئ�?��\�_?              �?                ��ۥ���?      �?       @      �?                       @               @       @       @                �#�d�Q�?��oHN�?                      �?        �z2~���?      �?       @                                       @       @       @              �?      �?��}�ɣ�?98ɛ���?      �?      �?      �?        H���@��?      �?                               @                                       @              @፿Po�?�C�j��?      �?              �?      �?�6��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �??�]�FR�?o�!��?                                              �?               @      �?      �?      �?      �?      �?      �?              �?      @�]�FR�?@}m[&?                                ��V��?      �?       @               @       @                                              �?      @I8O�)�?��P�U��?                      �?        �K=��?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?��N�Ա?��X�RR�?      �?              �?        �ԓ�ۥ�?              �?               @               @       @       @       @       @                z�rv��?���*���?      �?              �?        ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?�፿Po�?�$O��n?                                6��9�?      �?       @                               @                                      �?      @�%��}�?FP�۞��?                                F���@��?      �?       @      �?                                                              �?       @��Po��?��@7<�?      �?                                      �?              �?                                       @       @              �?       @8�B�]��?][L�̀?                                ��RO�o�?      �?              �?               @                               @              �?       @V�i���?�'�xV*�?                                              �?              �?                                                                       @q%�yO��?���F}�x?                      �?      �?$Zas �?      �?       @      �?                               @       @       @              �?      �?k1v��?϶�!��?                                F���@��?              �?                                                                      �?       @�p�Ȭ?�>�5��?      �?                                      �?              �?                                                              �?       @3NaJ̖�?Q^�}]x?                                �V�H�?      �?       @      �?                                       @       @                        �i����?�7J-�?      �?              �?      �?,l$Za�?      �?                               @               @                              �?        ]!ї�V�?޿R�ͯ�?                                �z2~���?      �?       @                                       @       @       @      �?              @��#�d��?����-9�?      �?                        �]�����?      �?       @      �?                               @       @       @      �?      �?       @.�jL��?m8�����?                                ��ۥ���?      �?       @      �?               @       @               @       @      �?      �?        Y7���?�x�4��?      �?              �?      �?Zas �
�?      �?              �?               @       @       @       @       @      �?              �?�� Q�E�?�	ܡ��?                      �?      �?H���@��?      �?       @                       @               @       @       @       @                ���Up�?����t��?                                �D+l$�?      �?       @               @                       @               @      �?                +�oM�?.�u���?                                �@�6�?              �?               @       @               @               @                      �?�������?�C���?      �?                        �D+l$�?      �?                                       @       @       @                      �?       @���Z��?j��q�r�?                                �@�6�?      �?       @      �?       @                                                      �?      �?���[�?��r¸l�?      �?                        F���@��?      �?       @      �?                                       @       @              �?       @=���&�?#�&f[)�?      �?              �?        Zas �
�?      �?              �?               @       @       @               @                      �?Q�E�*�?3?��?      �?              �?              �?      �?       @               @               @       @       @       @       @              �?��ds��?�Y��$o�?      �?                        [as �
�?              �?                               @               @       @      �?      �?       @yO�0@�?&{
�69�?      �?              �?        H���@��?      �?       @      �?               @                       @       @              �?        ��?y4��?�/׽~��?      �?              �?      �?��RO�o�?      �?              �?               @               @       @                      �?       @����_��?�Z#PB��?              �?      �?        !�
���?      �?       @      �?       @                                                      �?       @1�����?������?      �?              �?      �?p�z2~��?      �?              �?       @               @                       @                       @�^!ї��?{-�Fj�?                      �?        �V�H�?              �?               @       @                       @                               @O�0@�b�?����W.�?                      �?        ���V،?      �?                       @                                       @              �?      @e�����?��xI�?              �?      �?        ��RO�o�?      �?       @      �?                                       @       @      �?      �?      �?�>|]��?�K�]t�?      �?                        F���@��?      �?       @      �?                       @               @                      �?       @��ǰ2��?�Nʿ��?      �?              �?        3~�ԓ��?      �?       @      �?                               @                      �?      �?       @�I�:Bl�?��e=4�?                              �?ܥ���.�?              �?                       @       @                       @                      �?O�0@�b�?��@	��?      �?              �?      �?�'�K=�?      �?               @      �?      �?      �?      �?      �?      �?       @              @nC��x�?�k��O�?                                              �?              �?                                                                      @�/�����?�t�Y=�x?      �?                        H���@��?      �?                       @       @               @       @       @              �?      @T�n�W�?'w7���?              �?                ���V،?      �?              �?                                                                       @L�*g��?�z'y�?      �?                        ?���@��?      �?                               @                                                      @!�iŽ�?�Z��h�?                      �?      �?�
��V�?      �?               @      �?      �?      �?      �?      �?      �?       @              @Z��2�?�_- Q��?      �?      �?      �?        ��ۥ���?      �?                                       @       @                      �?              �?��7q��?%�5-N(�?                                ܥ���.�?      �?              �?               @                                      �?               @_W-��?�����?                                e�v�'��?      �?       @      �?               @       @       @       @       @                       @aѲ
n��?��C$�?      �?              �?        �ԓ�ۥ�?      �?       @      �?                       @               @       @      �?                �۴���? ���y1�?      �?              �?      �?3~�ԓ��?      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?t+�oM�?j=o��?      �?                        ��ۥ���?      �?       @               @       @       @       @               @       @                r�g�L��?�Ak�5�?                      �?        ?���@��?              �?               @                                                      �?       @
�X����?���V/�?                              �?�V�H�?      �?              �?       @       @               @       @       @      �?      �?        s[ݧ���?��KI��?                                6��9�?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����`�?ɞB�M��?                      �?        �]�����?      �?       @      �?               @                                                       @*L����?��_�p��?      �?                                      �?              �?                                               @                       @4�G�Ɉ�?0�ֺ�|?                                ���Vج?              �?                               @                       @                       @�w����?ݨǟn��?      �?      �?                F���@��?      �?       @      �?               @       @               @       @              �?       @]I`�:�?YC<����?                      �?        H���@��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�Y;���?31�J��?                      �?      �?P�o�z2�?      �?       @      �?                                       @              �?      �?       @	�M+��?�l����?                                �'�K=�?      �?              �?               @                                                       @:x��B�?�$�ć�?      �?              �?        ��.�d��?      �?                       @       @                       @       @      �?      �?      @/M��o2�?kI؀h�?                      �?      �?      �?      �?       @               @               @       @       @       @       @              �?��a�(�?������?              �?                [as �
�?      �?              �?       @                                                      �?      �?���G���?��;��?                      �?      �?�D+l$�?      �?       @      �?               @       @               @       @      �?      �?       @�g{���?�g<�?      �?                        !�
���?      �?       @      �?       @       @                       @              �?      �?       @����_�?��z:��?              �?                 �
���?      �?       @                                       @               @              �?       @MaJ̖p�?�9.�� �?      �?      �?      �?      �?�6��?      �?       @      �?               @                       @       @                       @�3i�ae�?�P��~�?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @F��1��?��ֺ�?      �?              �?      �?      �?      �?       @      �?       @       @               @               @       @      �?      �?�Wc"=P�?_���i��?      �?              �?      �?6���?      �?       @      �?                       @       @       @       @      �?      �?        )���G��?,�H��?                                �'�K=�?      �?                               @                                                       @�ti��|�?I\��5�?                                �]�����?      �?       @                       @       @       @       @       @      �?              �?�vAI�?����T��?                                F���@��?      �?                       @       @               @               @                        ��9���?�3&�GS�?      �?              �?      �?��ۥ���?      �?              �?       @       @       @       @       @       @       @              �?�MF���?�<|.b��?      �?      �?                ���V،?              �?                                                                      �?      @h#���?���qU!k?                                �V�H�?      �?                                                               @      �?              �?;�^!��?�0���?                      �?        �K=��?      �?       @               @       @       @                       @      �?              @��8j��?������?      �?                        H���@��?      �?       @      �?                                                              �?        ����9��?� W-V�?      �?              �?      �?F���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?        �����`�?��$�k�?      �?              �?      �?��V��?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?Y�)L�ْ?�q��Ʊ?                      �?      �?��V��?      �?       @               @       @               @       @       @       @      �?        jŽ�,u�?b���0�?                                ���V؜?      �?              �?                       @                                      �?      @F��s��?R��?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @���C�?ݘ<$3(?                              �?�z2~���?      �?       @      �?       @                                                      �?       @c=kg��?��x��M�?      �?                        �z2~���?      �?              �?       @               @               @       @      �?      �?      �?k1v��?'|�M%��?      �?                        �z2~���?      �?               @      �?      �?      �?      �?      �?      �?                       @9�%��}�?��eR�?      �?              �?      �?>�]���?      �?       @               @       @               @               @       @      �?      �?
n��W�?�֧�T�?      �?              �?      �?P�o�z2�?      �?              �?       @       @       @               @       @       @      �?      �?�w����?����?                      �?        3~�ԓ��?      �?       @      �?               @       @               @       @      �?      �?       @���-�j�?�eP�?      �?                                      �?              �?               @                               @              �?       @�_���@�?lߤJ?      �?              �?      �?H���@��?      �?       @      �?                                       @                               @�s��2�?�K¥�H�?      �?              �?        ��RO�o�?      �?                               @               @                              �?       @�G�Ɉ��?{A�;@�?                      �?        �
��V�?      �?       @      �?       @                               @                      �?        �hY7��?
��2�>�?                                {2~�ԓ�?              �?               @                       @       @       @      �?      �?        �
n���?0t];`�?      �?                      �?�z2~���?      �?       @      �?                                                              �?      �?*g���?<p�۹/�?      �?              �?      �?��ۥ���?      �?                               @               @       @       @       @      �?      �?����U��?�.'����?      �?                        F���@��?      �?       @      �?                                       @       @              �?       @m��W�?��{i�8�?                      �?      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?                �%��}�?y�V�7�?                                6��9�?      �?       @               @       @       @       @       @                      �?      �?��䶺O�?>�)���?      �?              �?                      �?              �?                                       @                      �?       @��r�9��?@f3­/}?      �?      �?      �?        $Zas �?      �?       @      �?               @       @               @       @              �?       @O|x�/��?�N+OT��?                      �?      �?3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?��N�ԑ?�7B�X��?                                ��.�d��?              �?               @       @               @                       @              @R�&#��?A:�F���?              �?                3~�ԓ��?      �?                               @               @                                        �5A .�?�Yԭ���?      �?                                      �?              �?                               @                              �?      @j�����??ښo;z?      �?                                      �?               @      �?      �?      �?      �?      �?      �?                      @��%��}z? �<$3�>      �?                      �?	��V��?      �?                       @                                                      �?      @ e��h�?��q��u�?                      �?      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                n��W�?jՓ��?      �?                        (�K=�?      �?       @      �?       @                       @       @       @       @      �?      �?'Y��M�?q��ҳ�?      �?                              �?              �?               @       @       @       @       @       @       @      �?        ��g{��?��<��j�?              �?                              �?              �?                                                              �?       @��6���?l�O7WKx?                      �?        �D+l$�?      �?              �?               @               @       @       @       @      �?      @��_���?�:7�6�?                      �?      �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?       @              @�፿Po�?��5�.��?                                �o�z2~�?      �?       @      �?                                       @       @      �?      �?        ��1��?�x��0�?                      �?        �K=��?      �?               @      �?      �?      �?      �?      �?      �?       @              @�U�����?��4�q�?                                ��.�d��?      �?                       @               @       @                      �?              �?\�yjH�?��3�'T�?                      �?      �?(�K=�?      �?       @      �?       @       @       @       @       @       @       @      �?      �?��a/�?��a���?                                ��RO�o�?      �?                                               @               @      �?              �?i1v��?M ��rF�?                      �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @      �?      �?�J���?�^�IJ��?      �?              �?      �??���@��?              �?               @                               @                              �?�E�X���?��eI9�?      �?                        	��V��?      �?               @      �?      �?      �?      �?      �?      �?       @              �?����'t�?U{��?                                �
��V�?      �?                                                                      �?                �?����C�?      �?                      �??���@��?      �?       @      �?                               @                                      �?�:]���?�	�7釢?              �?      �?        v�'�K�?      �?       @                       @       @               @       @       @      �?        ��r�9��?�J~X_�?      �?              �?      �?ܥ���.�?      �?       @      �?       @       @       @       @       @       @       @              �?�}��?`v.!�?      �?              �?              �?      �?                       @       @       @       @       @       @       @              @#���?pfC�V5�?      �?                      �?���V،?      �?       @               @       @                                                        ��8�)1�?��K�]�?      �?                        p�z2~��?      �?              �?                               @       @       @              �?       @4�돗��?]��Y�?      �?              �?        e�v�'��?      �?                       @       @                       @       @       @      �?        9ֳv&��?,W���?      �?              �?      �?      �?              �?               @       @       @       @       @       @       @      �?      �?UH�%���?�t2||�?      �?              �?        Zas �
�?      �?       @      �?                                                              �?       @/M��o2�?ύ^�IJ�?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @      �?      �?        ���,���?      �?                      �?        !�
���?      �?       @      �?                       @               @       @      �?      �?       @��l	��?�� *3�?                                6��9�?      �?                               @                       @              �?               @��	�p�?c��?tR�?                                ��ۥ���?      �?       @               @                                              �?              @�ߚ ��?��2K���?                                H���@��?      �?       @      �?               @                       @       @              �?       @��2�?PB���~�?                      �?        (�K=�?              �?                       @       @       @       @       @       @                ��B�/�?7YBq/��?                                ���V،?      �?                                                                              �?      @)g��1�?���V/z?      �?                        3~�ԓ��?      �?               @      �?      �?      �?      �?      �?      �?      �?              @-h#���?	2�e�?                      �?      �?��Vؼ?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����`�?�I,��$�?                                �ԓ�ۥ�?      �?       @      �?                               @       @       @              �?        䛌8j��?�<����?      �?              �?        !�
���?      �?       @      �?       @       @                               @      �?      �?      �?M��o2��?�>�5��?      �?                        �]�����?              �?                               @       @               @      �?               @���"X~�?ԈDX�?�?      �?      �?      �?        Zas �
�?      �?              �?                       @       @               @              �?       @^!ї�V�?���+x�?      �?              �?      �?��ۥ���?      �?       @               @       @       @       @       @       @       @               @����?�tX�I�?      �?                        ���V؜?      �?                                               @                              �?      @�����`�?�RH���?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?                      @��N�ԑ?��N��?                      �?      �?H���@��?      �?                       @               @       @                                        6&����?�0��1�?      �?                        �V�H�?      �?       @      �?               @       @               @              �?      �?      �?p2��g�?w�"BC�?      �?                      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @                F��1��?�9��%��?                      �?      �?p�z2~��?      �?                               @               @               @       @                �;x��?�K���?                                �@�6�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�X����?�	4Lo�?      �?                                      �?                                                                              �?       @�Y e�?��$�f?      �?                        �V�H�?      �?       @      �?                                                                        �<�^�?A8}���?      �?              �?      �?[as �
�?      �?       @      �?       @               @               @              �?                t J�h�?Ƀ��?      �?                                              �?                                                                      �?       @qi��|��?G,˽H?      �?      �?                �ԓ�ۥ�?      �?       @      �?                                       @       @              �?       @��f��?��,���?      �?                      �?��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @��*��?�֔LO)�?      �?                        ���Vج?              �?                       @                       @       @              �?      @w�����?Hm\2��?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?                       @F��1��?�1� �r?      �?              �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @                h#���?CmA��H�?                              �?6��9�?      �?       @               @               @       @               @      �?              �?���G���?������?      �?                      �?              �?       @                                                                      �?       @yO�0@�?C�{�m�m?      �?              �?      �??���@��?      �?              �?                                                              �?      @���U�?��~�rq�?      �?                        ���V؜?      �?       @                                                                                +���?y�?߈�(��?              �?      �?        ���@��?      �?       @      �?                               @       @       @      �?      �?       @H���<�?ҫS��?      �?              �?        p�z2~��?      �?               @      �?      �?      �?      �?      �?      �?      �?                �d�Q�ϐ?g�cV�L�?                      �?        �ԓ�ۥ�?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�?�t�\�?              �?      �?      �?�z2~���?              �?                                       @                              �?      @�S��%�?������?                                ���V؜?      �?               @      �?      �?      �?      �?      �?      �?              �?      @��N�ԑ?�Q��Ft?      �?                        6���?      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?h#���?F͙(�?                                p�z2~��?      �?              �?       @                                                              �?���6�?p�k��
�?                      �?        �@�6�?      �?              �?                               @       @                      �?       @�����?���.���?      �?              �?        �ԓ�ۥ�?      �?                                                                              �?        ��J��?R%�*&"�?                      �?      �?�z2~���?      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�U�����?��2H��?      �?                      �?��V��?      �?       @      �?       @               @                       @              �?        �������?F�^z�?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?      �?                Y�)L�ْ?5��r�?                                p�z2~��?      �?       @      �?                       @               @                      �?      �?�����?]���lV�?                                ���V؜?      �?                               @               @       @       @              �?       @���H*�?P���B��?      �?                                      �?                                               @                                      @��*��?K+� n�l?              �?                �]�����?              �?               @       @                                              �?      �?����[�?�����?                      �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ]����`�?��L$ �?                      �?        F���@��?      �?              �?                                       @                      �?       @����?���L�z�?                                �]�����?      �?                               @       @               @              �?                ��M+��?�5ݪ�?      �?                                      �?                                                                              �?      @��g{�?	�6�mi?                      �?      �?6��9�?      �?       @      �?               @                       @                      �?       @r�9ֳv�?-5���?      �?                        �@�6�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @8�]�FR�?;`���}�?                      �?        ��ۥ���?      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�U�����?ap9#{k�?                                	��V��?      �?               @      �?      �?      �?      �?      �?      �?                      �?^��Z��?\��e��?                                v�'�K�?              �?               @       @       @       @                       @      �?      @����,��?_ɮ8cS�?                              �?�ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?                ����[�?�/��3��?                      �?      �?              �?               @      �?      �?      �?      �?      �?      �?                      @n��W�?�^/��"?                                ���Vج?      �?                       @                       @       @                      �?       @w�D_r[�?��M�n��?      �?              �?        �ԓ�ۥ�?      �?       @      �?                               @               @              �?        t3NaJ��?P�r5�?                                ���V؜?      �?              �?       @                                                      �?       @9ֳv&��?Qn�&c�?              �?                ?���@��?      �?       @      �?                       @                       @              �?       @5\.2�z�?7�����?      �?              �?      �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?       @                �c=kgҮ?����d��?      �?                        e�v�'��?      �?       @               @               @       @       @       @       @                ����!��?`H�mj�?              �?                ��RO�o�?      �?              �?       @       @                                                       @���Z�K�?��Q}G�?                      �?        (�K=�?              �?               @               @       @               @       @      �?        h#���?��|!.��?      �?                        p�z2~��?      �?                       @                                                      �?        B�/����?׬�̱��?                      �?      �?�z2~���?      �?       @      �?                                               @                       @����q�?�x���Q�?      �?      �?                ?���@��?      �?              �?                                                                       @�vAIE�?��w$��?      �?              �?        ���V؜?              �?                                                       @              �?       @w�Τ=��?}��m!�?                      �?        �K=��?      �?                                               @                                        :�X�?~�gj��?                      �?      �?�RO�o��?      �?                               @       @       @       @       @       @      �?        r�g�L��?ySm\2�?      �?                                      �?              �?               @                                              �?       @,�����?��c|Az?                                ���V؜?      �?              �?               @                       @       @              �?       @{]�;x�?H���?      �?              �?      �?F���@��?              �?               @       @       @               @       @                      @�E�X���? =LLg�?                      �?        �ԓ�ۥ�?      �?                                               @                              �?      @ e��h�?-���.J�?              �?                �ԓ�ۥ�?      �?       @      �?               @               @                              �?       @b�(Ţe�?Ѻ����?                                H���@��?              �?                               @       @       @       @      �?               @�
����?'��%��?      �?              �?      �?      �?      �?       @      �?       @       @       @       @               @       @      �?      �?ߚ ���?�����{�?      �?                        ?���@��?      �?                       @               @                                               @ƽ�,u��?����?      �?                        !�
���?      �?               @      �?      �?      �?      �?      �?      �?      �?               @�]�FR�?�iy�=7�?      �?              �?        ��V��?      �?       @      �?       @       @       @                              �?               @�d�#��?#e�S@<�?                                              �?       @      �?               @                       @       @              �?      �?��2�?v͑�?�?      �?                        v�'�K�?      �?       @      �?               @               @       @       @      �?      �?       @�N��b�? 8]ϓC�?                      �?      �?!�
���?              �?                               @       @       @       @      �?      �?       @z����"�?��TN;E�?                      �?      �?�V�H�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?�፿Po�?}�AĿ�?                                �ԓ�ۥ�?      �?       @               @               @       @       @       @       @      �?      �?��>|]�?�m	���?                                	��V��?      �?              �?               @                       @                      �?       @kg����?<���Z�?      �?                        �
��V�?      �?              �?       @       @                       @       @      �?      �?      @�=�� Q�?4�ߺ�n�?                                ���Vج?      �?               @      �?      �?      �?      �?      �?      �?                      @����[�?\Z ��n�?                      �?      �?�K=��?      �?               @      �?      �?      �?      �?      �?      �?                      @����'t�?\�a����?      �?              �?        �ԓ�ۥ�?      �?                       @       @       @                                              @Xc"=P9�?."Ӵ�0�?                                p�z2~��?      �?       @      �?                               @               @              �?       @�r�9ֳ�?�I�����?      �?              �?      �?p�z2~��?      �?                       @       @               @               @              �?      �?p�l�?�؞]��?      �?              �?      �?6��9�?      �?               @      �?      �?      �?      �?      �?      �?       @              @#w\I`ޓ?�ϖǥ?              �?                ���Vج?      �?              �?       @       @                                                       @�AQ�s��?M7��r�?                                ���V،?      �?               @      �?      �?      �?      �?      �?      �?              �?        �Y;���?�^�)�c?                      �?      �?���@��?      �?       @                       @       @       @       @       @      �?      �?      �?��Kn���?�[�C���?      �?              �?      �?�'�K=�?      �?                       @                                                      �?      �?����?F�r5�?      �?              �?      �?P�o�z2�?      �?       @       @      �?      �?      �?      �?      �?      �?       @                ���6�?�p�j<��?      �?                        F���@��?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�U����|?�P~~�h�?                      �?      �?v�'�K�?      �?                                               @                      �?      �?      �?��r�9��?���Fm��?      �?                        �K=��?      �?                               @                                              �?       @፿Po�?�D]KV�?                                6��9�?      �?       @      �?       @       @                               @              �?       @?(�tN|�?���As&�?      �?                                      �?                                                                              �?        z+�oM�?����
�g?      �?              �?              �?      �?       @      �?       @       @       @       @       @       @       @              �?s����?�=71��?                      �?      �?      �?      �?                       @       @       @                       @       @              �?����`�?����?      �?              �?      �?(�K=�?      �?       @                       @       @       @       @       @       @      �?      �?l�\d��?�=�@���?                                ���V،?      �?              �?                                                                       @3NaJ̖�?� �'w�?      �?              �?        (�K=�?      �?       @               @               @       @               @       @              �?%fK8O��?t}'�;�?      �?                        ��Vؼ?      �?       @      �?                                                              �?       @#�6��w�?\������?                                ��ۥ���?      �?               @      �?      �?      �?      �?      �?      �?      �?              @�%��}�?f�4ȱ?      �?                        	��V��?      �?                       @       @                                      �?              @�%��}�?4�{Ck�?                      �?      �?���.�d�?      �?       @      �?       @       @       @       @       @       @      �?               @�u�4�G�?�Z3F��?      �?                        ��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?nC��x�?��&(z�?              �?      �?                      �?                                                                                       @*g���?�ppTV�i?      �?      �?      �?        F���@��?      �?       @      �?                                       @       @              �?        IE����?�� @�z�?      �?                        P�o�z2�?      �?       @      �?       @       @       @       @       @       @      �?      �?      �?`r[ݧ��?5m&̣��?      �?                      �?��RO�o�?      �?               @      �?      �?      �?      �?      �?      �?       @              �?^��Z��?�QI���?      �?      �?      �?        �@�6�?      �?              �?               @                               @              �?       @T�@ʾ��?V�_����?                      �?        ��V��?      �?                       @               @                                      �?      @�a/��?4P����?              �?      �?        [as �
�?              �?               @       @       @                       @      �?      �?      �?+���?y�?~����?                                              �?              �?                                       @                      �?       @!�iŽ�?Z�a}?                      �?      �?e�v�'��?      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        ��w����?p�a�ދ�?                      �?        ���Vج?      �?              �?                                                              �?       @� �;�$�?`
��?                      �?        ?���@��?      �?       @      �?               @                       @                      �?       @嶺O_�?�2�fFz�?      �?              �?        (�K=�?      �?       @               @                       @       @       @       @      �?      �?�ڙ�ǰ�?^��ձv�?      �?                        �@�6�?      �?              �?                               @                              �?       @��N���?�N>���?              �?                �ԓ�ۥ�?      �?               @      �?      �?      �?      �?      �?      �?      �?                E�(Ţe�?"�y�̹�?      �?                        Zas �
�?      �?               @      �?      �?      �?      �?      �?      �?              �?      @^��Z��?�2@g�?                      �?              �?              �?               @       @       @       @       @       @       @                ��@���?��F}��?                      �?      �?Zas �
�?      �?       @      �?       @       @       @       @       @       @       @              �?Z.2�z��?ʑ��?�?       �t�b�n_samples_fit_�M:�_tree�N�_sklearn_version��1.2.2�ub.