��       �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�K*�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�
customerID��gender��SeniorCitizen��Partner��
Dependents��tenure��PhoneService��MultipleLines��InternetService��OnlineSecurity��OnlineBackup��DeviceProtection��TechSupport��StreamingTV��StreamingMovies��Contract��PaperlessBilling��PaymentMethod��MonthlyCharges��TotalCharges�et�b�n_features_in_�K�
n_outputs_�K�classes_�hhK ��h��R�(KK��h �i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���hEC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��hE�C       �t�bK��R�}�(h	K�
node_count�M��nodes�hhK ��h��R�(KM���h �V56�����R�(Kh$N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hghEK ��hhhEK��hihEK��hjh �f8�����R�(KhFNNNJ����J����K t�bK��hkhuK ��hlhEK(��hmhuK0��uK8KKt�b�B��        �                   �?���%���?           �@       3      	             �?n��"O�?           �@                       ����?H6�(���?0           `�@       �                    �?~��6��?�           ��@       �                 �|�?XK�~���?�           py@       q                 �Ӻ}?�j4����?R            u@       T                 �Ӻm?l��@���?�             e@       S                    �?��|��L�?s            �\@	       J                    �?���
��?k            �Z@
       G                    �?      �?^            �W@       D       
             �?v ��?V            �U@       /                 `��?     ��?P             T@       ,                    �?�q���?0             H@                           L�@���Q��?(             D@                           H�@���y4F�?             3@                           �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @                        �J�g?      �?             0@                           �@z�G�z�?
             $@������������������������       �                     @                           ɡ@���Q��?             @                        �� �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                        ��DE?և���X�?             5@������������������������       �                      @       #                   �?p�ݯ��?             3@                            y�@      �?              @������������������������       �                     @!       "                 �(�?�q�q�?             @������������������������       �                      @������������������������       �                     �?$       %                 �
n�?�eP*L��?             &@������������������������       �                     @&       +                    ��@      �?              @'       *                    �?����X�?             @(       )                    4�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?-       .                 ����?      �?              @������������������������       �                     @������������������������       �                     �?0       A                    �?     ��?              @@1       <                 @5�?�<ݚ�?             ;@2       ;                    N�@��2(&�?             6@3       4                    1�@�����?             5@������������������������       �                     (@5       6                    ��@�<ݚ�?	             "@������������������������       �                     �?7       :                 �F�?      �?              @8       9                  �=�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?=       @                    �?���Q��?             @>       ?                    ^�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @B       C                   �ɳ@z�G�z�?             @������������������������       �                     @������������������������       �                     �?E       F                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @H       I                   �+�@      �?              @������������������������       �                     @������������������������       �                     �?K       R                    �@8�Z$���?             *@L       Q                   ��@����X�?             @M       N                 p@��?r�q��?             @������������������������       �                     @O       P                 0��h?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @U       h                 @؋�?������?6             K@V       W                    h~@��r._�?)            �D@������������������������       �                     �?X       g                    ��@R���Q�?(             D@Y       b                    �?�ݜ�?'            �C@Z       [                  &�t?l��\��?"             A@������������������������       �                     5@\       a                   ���@�θ�?             *@]       ^                 �� �?�C��2(�?             &@������������������������       �                      @_       `                    ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @c       d                 ���?���Q��?             @������������������������       �                      @e       f                 `��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?i       j                  ��?��
ц��?             *@������������������������       �                     @k       p                 ��!�?�q�q�?	             "@l       m                    �?؇���X�?             @������������������������       �                     @n       o                 @�-s?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @r       �                 ��8�?|ƀQK��?�             e@s       �                    �?X�<ݚ�?�            @d@t       �                    x�@���A��?�            �a@u       �                  ���?z�G���?P             T@v       �                 ����?�eP*L��?B            �P@w       ~                    �?X�Cc�?             <@x       }                    �@     ��?             0@y       |                 ���?�r����?             .@z       {                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?       �                 `h�?�q�q�?             (@�       �                    �?�z�G��?
             $@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   J�?�����?&             C@������������������������       �                     @�       �                 ��f�?���|���?!            �@@������������������������       �                      @�       �                    ��@�4�����?             ?@�       �                    B�@D�n�3�?             3@�       �                  C1�?     ��?             0@�       �                 P��?�eP*L��?             &@�       �                 @��?�q�q�?	             "@�       �                 xǡ?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?r�q��?             (@������������������������       �        
             $@������������������������       �                      @�       �                    �?d}h���?             ,@������������������������       �                      @�       �                    j�@�8��8��?             (@������������������������       �        	             "@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �@�4�����?>             O@�       �                 �̱�?z�G�z�?             >@������������������������       �                     �?�       �                   �t�@д>��C�?             =@������������������������       �                      @�       �                 �C��?���N8�?             5@�       �                 �0@�?z�G�z�?             4@�       �                 ���?�q�q�?             (@�       �                    �?z�G�z�?
             $@�       �                    �?�����H�?	             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �a�@     ��?              @@������������������������       �                     @�       �                    �?�q�q�?             ;@�       �                    �?�GN�z�?             6@�       �                  ���?�t����?             1@�       �                   �[�@      �?             0@�       �                 ���?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     �?�       �                    �?���Q��?             @�       �                 @��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                 �ї?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    ��@��Q��?             4@�       �                 ����?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?؇���X�?             ,@�       �                    �?$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?������������������������       �                     @�       �                 P�c�?&�a2o��?E            @Q@�       �                 p���?d�;lr�??            �O@�       �       
             �?�d�����?&             C@�       �                    �?��}*_��?             ;@�       �                 ��8�?�q�q�?             8@�       �                  �Ǩ?�8��8��?             (@������������������������       �        
             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             (@�       �                 ��a�?����X�?             @������������������������       �                     �?�       �                 �v�?r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@�       �                    @`2U0*��?             9@������������������������       �                     4@�       �                 �-��?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       1                ���?䖏��J�?]           �@�       �                 `p�?ԳC��2�?�             f@������������������������       �                     ?@�                       ��Dz?д>��C�?�             b@�                         ���@�E��ӭ�?6             K@�       �                    �?�MI8d�?%            �B@������������������������       �                     �?�       �                    �K@4?,R��?$             B@������������������������       �                     �?�       �                    (�@(N:!���?#            �A@������������������������       �                     *@�       �                    4�@"pc�
�?             6@������������������������       �                     �?�       �                 �'t�?؇���X�?             5@�       �                    ��@      �?              @������������������������       �                     �?������������������������       �                     �?�                        p@��?�KM�]�?             3@������������������������       �                     (@                         �?����X�?             @                        �5�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                        ���@��.k���?             1@                      $3x?�q�q�?             (@������������������������       �                     �?	                       v>z?���!pc�?             &@
                         �?z�G�z�?
             $@                         @���Q��?             @                       ֘�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?                      P���?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                          ,�@L�[2[
�?[            �V@                         ̌@      �?             8@������������������������       �        
             $@                      �h��?և���X�?             ,@                         �?�q�q�?             (@                         �?z�G�z�?
             $@������������������������       �                     @                         �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @!      &                �/��?�L#���?C            �P@"      #                   �?P�Lt�<�?&             C@������������������������       �                      @@$      %                   S�@r�q��?             @������������������������       �                     �?������������������������       �                     @'      (                ��>}?ܷ��?��?             =@������������������������       �                     �?)      0                �ߵ�?@4և���?             <@*      /                �(��?�r����?             .@+      .                   �?@4և���?             ,@,      -                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             "@������������������������       �                     �?������������������������       �                     *@2      �                � Q�?"�{	�?�           �z@3      p                  �ϲ@X)0���?�            �`@4      E                   �?�ހ��?^            �W@5      @                 KS�?�GN�z�?             6@6      =      
             �?�t����?             1@7      8                   �?��S�ۿ?             .@������������������������       �        
             $@9      :                 �Ҏ?z�G�z�?             @������������������������       �                     @;      <                XUU�?      �?              @������������������������       �                     �?������������������������       �                     �?>      ?                   �?      �?              @������������������������       �                     �?������������������������       �                     �?A      D                   ��@���Q��?             @B      C                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @F      o                P�@�?)O���?H             R@G      n                �@�?��z4���?E            @Q@H      a                   x�@������??            �O@I      J                �'�?�+��<��?+            �E@������������������������       �                     @K      V                   Ɯ@��+��?%            �B@L      M                p���?���|���?             6@������������������������       �                     @N      O                �yO�?��S���?             .@������������������������       �                      @P      Q                }�?�n_Y�K�?             *@������������������������       �                     @R      S                �}��?      �?              @������������������������       �                     @T      U                �8��?���Q��?             @������������������������       �                      @������������������������       �                     @W      \                0#��?�q�q�?             .@X      [                   c�@      �?              @Y      Z                   4�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @]      `                   �?և���X�?             @^      _                0'+�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @b      m      
             �?��Q��?             4@c      l                �-&�?�E��ӭ�?             2@d      k                ��0�?������?             1@e      f                �,�?���Q��?
             $@������������������������       �                     @g      h                p.	�?և���X�?             @������������������������       �                     @i      j                �!�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @q      �                �8��?���Q��?(             D@r      s                �P��?\X��t�?             7@������������������������       �                     @t      {                   �?�����?             3@u      z                0�)�?      �?
             $@v      w                   �?      �?              @������������������������       �                     @x      y                ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @|                         �?�����H�?	             "@}      ~                   Ѷ@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                ��޶?@�0�!��?             1@�      �                   �?      �?             0@������������������������       �                     (@�      �                ���?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�      �                   �?���v{�?'           pr@�      �                 J��?���W�?�            �a@�      �                   @�>����?             ;@�      �                Pn��? �q�q�?             8@�      �                �=��?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     1@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                � W�?�û��|�?s            �\@�      �                p��?"pc�
�?             &@������������������������       �                      @������������������������       �        	             "@�      �                  ��@$��m��?h             Z@�      �                  �#�@�y�ʍ+�?\             W@�      �                ��?8�$�>�?V            �U@�      �                 s�?�D��?1            �H@�      �                �Y �?\X��t�?             7@�      �                  ���@�θ�?             *@�      �                   @ףp=
�?
             $@������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?�z�G��?
             $@������������������������       �                     @�      �                ���?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   �?ȵHPS!�?             :@������������������������       �                     3@�      �                   �?և���X�?             @�      �      
             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                ����?��%��?%            �B@������������������������       �                     @�      �                   d�@      �?              @@�      �                ����?ףp=
�?
             $@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                 |��?      �?             6@������������������������       �                     @�      �                `;��?D�n�3�?             3@�      �                   �?�<ݚ�?	             "@������������������������       �                      @������������������������       �                     @�      �                   �?���Q��?
             $@�      �                `p�?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                @���?r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�      �                 ���?��k����?�             c@������������������������       �                     @�                        �ƺ@�7�QJW�?�            �b@�                      �<�?ZՏ�m|�?�            `b@�                      ��ɸ?�@i����?�            @b@�      �                   �?��2(&�?�            �`@�      �                   �?�����?D             Q@�      �                  �Y�@8^s]e�?             =@�      �                   ذ@���Q��?             4@�      �                   ~�@      �?             0@�      �                   �?      �?              @�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                а2�?�����H�?	             "@�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   �?��-�=��?'            �C@�      �                ��6�?����X�?             @�      �                �v�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   �?      �?              @@�      �                   }�@XB���?             =@������������������������       �                     6@�      �      
             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                �Q��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                ��e�?     p�?@             P@������������������������       �                     9@�      �                пk�?�ݜ�?'            �C@������������������������       �                     �?�      �                   ��@�KM�]�?&             C@������������������������       �                     2@�      �                   �?z�G�z�?             4@�      �                �q�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                 4��?�t����?             1@�      �                ��s�?      �?              @������������������������       �                     �?������������������������       �                     �?�                          ��@��S�ۿ?             .@�      �                   %�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@                         �?X�Cc�?             ,@                      ��8�?      �?             (@������������������������       �                     �?            
             �?"pc�
�?             &@������������������������       �                     @                         ښ@      �?             @������������������������       �                     �?	      
                �C��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?                         '�@�q�q�?             @������������������������       �                      @������������������������       �                     �?      �                   �?�Wu�1��?<           �@      K                   �?Z'8of�?           `q@                      p�ҡ?���;�?r            �\@������������������������       �                      @                      ��?���X��?p             \@                         �?�����H�?             ;@                      ���?�z�G��?
             $@                       �1�?���Q��?             @                      � �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     1@      B                   �?ҳ�wY;�?U            @U@       1                   ��@և���X�??            �O@!      *                   ��@:ɨ��?!            �@@"      '                   ��@��
ц��?             *@#      $                   �?����X�?             @������������������������       �                     @%      &                   H�@�q�q�?             @������������������������       �                      @������������������������       �                     �?(      )                �!�?r�q��?             @������������������������       �                     @������������������������       �                     �?+      .                ����?R���Q�?             4@,      -                   �?��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@/      0                p��?���Q��?             @������������������������       �                      @������������������������       �                     @2      3                   ̭@*;L]n�?             >@������������������������       �                     @4      =                 �~�?�q�����?             9@5      <                   @X�Cc�?             ,@6      7                   �?      �?             (@������������������������       �                     @8      9                   �?      �?             @������������������������       �                      @:      ;                   @�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @>      ?                �Ű�?���!pc�?             &@������������������������       �                     @@      A                `_x�?���Q��?             @������������������������       �                     @������������������������       �                      @C      D                   \�@��2(&�?             6@������������������������       �                     �?E      F                   �?�����?             5@������������������������       �                     .@G      H                   �?�q�q�?             @������������������������       �                     @I      J                0O�?�q�q�?             @������������������������       �                      @������������������������       �                     �?L      m                 �q�?�p ��?�            �d@M      \                p��?�G�5��?E            @Q@N      S                �'��?4?,R��?$             B@O      P                ����?���Q��?             @������������������������       �                      @Q      R                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?T      U                   �?`Jj��?             ?@������������������������       �                     2@V      W                �`�?8�Z$���?             *@������������������������       �                     �?X      [                 �q�?�8��8��?             (@Y      Z                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             $@]      j                   ��@���|���?!            �@@^      i                @X��?      �?             8@_      d                ���?ҳ�wY;�?             1@`      a                   �?ףp=
�?
             $@������������������������       �                      @b      c                   �?      �?              @������������������������       �                     �?������������������������       �                     �?e      f                   �?����X�?             @������������������������       �                     �?g      h                   ��@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @k      l                p��?�q�q�?	             "@������������������������       �                     @������������������������       �                     @n      u                ����?�:nR&y�?_            �W@o      p                   �?      �?@             P@������������������������       �        /            �G@q      r                   w�@�t����?             1@������������������������       �                     ,@s      t                p�#�?�q�q�?             @������������������������       �                      @������������������������       �                     �?v      �                   '�@�חF�P�?             ?@w      x                �P�?�r����?             >@������������������������       �        
             $@y      ~                @lv�?z�G�z�?             4@z      {                   �?      �?             @������������������������       �                      @|      }                   �?      �?             @������������������������       �                     @������������������������       �                     �?      �                   �@@4և���?             ,@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?�                         �?�ʱOY��?&           0�@�      �                ����?�2l����?+           �r@�      �                   �?��#����?�            @l@�      �                �8��?dy�����?�            `c@�      �                ��8�?4�M�f��?f            �Y@�      �                0��?�q�q�?T             U@�      �                �AQ�?�������?D             Q@�      �                `��?b�2�tk�?6             K@�      �                @؀�?�z�G��?
             $@������������������������       �                     @������������������������       �                     @�      �                �N�?�X����?,             F@�      �                ���?|��?���?             ;@�      �                   �?      �?              @������������������������       �                     @�      �                �k��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                 �q�?p�ݯ��?             3@�      �                ����?�q�q�?             (@�      �                  �X�@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?�IєX�?             1@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@�      �                   X�@؇���X�?             ,@������������������������       �                     �?�      �                   �?$�q-�?             *@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�      �      
             �?      �?             0@������������������������       �                     &@�      �                `�+�?���Q��?             @������������������������       �                     @������������������������       �                      @�      �                  ���@�<ݚ�?             2@������������������������       �                     *@�      �                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                   �@�T`�[k�?5            �J@�      �                 ��?      �?              @������������������������       �                     @�      �                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                  �+�@:	��ʵ�?-            �F@�      �                   �?�����H�?$             B@�      �                p���?���!pc�?             &@�      �                P��?�����H�?	             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                �V�?`2U0*��?             9@�      �                ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     5@�      �                   �?X�<ݚ�?	             "@�      �                  �P�@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   ��@�ˡ�5��?G            �Q@�      �                �#��?�t����?3            �I@�      �                ���?�>4և��?             <@�      �                @���?H%u��?             9@������������������������       �                     *@�      �                0�v�?      �?             (@������������������������       �                     �?�      �                ����?"pc�
�?             &@������������������������       �                     �?�      �                  ���@ףp=
�?
             $@������������������������       �                     @�      �                   :�@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                Б��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                p�?�nkK�?             7@�      �                ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@�      �                   ��@�z�G��?             4@�      �                   �?      �?
             $@�      �                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                @�c�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                ���?ףp=
�?
             $@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                   �?��-*��?I            @R@�      �      
             �?�LQ�1	�?             7@�      �                �}��?      �?              @������������������������       �                     @�      �                   ��@���Q��?             @�      �                P��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                   �?z�G�z�?             .@�      �                ���?      �?              @������������������������       �                     @�      �                 �E�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                       ����?���Q��?2             I@                         �?r�q��?             (@������������������������       �                     �?                         �?�C��2(�?             &@������������������������       �        	             "@                      ���?      �?              @������������������������       �                     �?������������������������       �                     �?      	                 ��?�\��N��?&             C@������������������������       �                     @
                         R�@����e��?!            �@@������������������������       �                     @                      Pm?�?|��?���?             ;@                      �Jk�?�	j*D�?             *@                      �<�?      �?             @������������������������       �                     @������������������������       �                     �?                       ���?�����H�?	             "@������������������������       �                     @                         f�@      �?              @������������������������       �                     �?������������������������       �                     �?                      @q�?����X�?             ,@                      `(��?ףp=
�?
             $@������������������������       �                     �?������������������������       �        	             "@                         d�@      �?             @������������������������       �                     @������������������������       �                     �?      P                   �?Hث3���?�           �@      /                   �?�q�q�?T             U@      ,                   
�@���@��?%            �B@       !                @w\�?��Q��?             4@������������������������       �                      @"      #                �1��?�E��ӭ�?             2@������������������������       �                     @$      '                �~�?�eP*L��?             &@%      &                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @(      +                �3��?r�q��?             @)      *      
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @-      .                hM�?�IєX�?             1@������������������������       �                     �?������������������������       �                     0@0      A                   �?�[�IJ�?/            �G@1      <                   Q�@�q�q�?             8@2      ;                ����?�<ݚ�?             2@3      8                   �?@�0�!��?             1@4      7                   ��@$�q-�?             *@5      6                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@9      :                   ڪ@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?=      >                �8��?�q�q�?             @������������������������       �                     @?      @                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?B      C                ��>�?
;&����?             7@������������������������       �                     @D      E                @ �?�G�z��?             4@������������������������       �                     @F      K                   >�@     ��?             0@G      H                   �?      �?              @������������������������       �                     @I      J                ����?      �?             @������������������������       �                      @������������������������       �                      @L      M                   �?      �?              @������������������������       �                     @N      O                   �?      �?             @������������������������       �                     �?������������������������       �                     @Q      �                PUU�?� ��	��?�           pz@R      a                �ڽ?p�v>��?^            �W@S      T                `K�?�q�q�?             8@������������������������       �                     @U      V                   ܕ@�q�q�?             5@������������������������       �                     @W      X                   ��@     ��?             0@������������������������       �                      @Y      ^                   �?X�Cc�?             ,@Z      [                ��=�?z�G�z�?
             $@������������������������       �                     @\      ]                ����?      �?             @������������������������       �                      @������������������������       �                      @_      `                   �?      �?             @������������������������       �                     @������������������������       �                     �?b      g                �N.�?z�G�z�?F            �Q@c      f                @q��?(;L]n�?             >@d      e                4��?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@h      i                �^�?�G�z�?(             D@������������������������       �                     @j      {                @�5�?����>�?%            �B@k      r                Ц�?�û��|�?             7@l      m                   T�@"pc�
�?             &@������������������������       �                     �?n      q                 ���?ףp=
�?
             $@o      p                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @s      x                P���?�q�q�?             (@t      w                   �?؇���X�?             @u      v                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @y      z                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?|      }                   q�@@4և���?             ,@������������������������       �                     &@~                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      $                �q�?�^�Q��?I           �t@�      �                   ^�@�����?+           �r@�      �                   ��@ؓ��M{�?n            �[@�      �                ��?�xGZ���?i            @Z@�      �                   �_@���/��?O            �S@������������������������       �                     @�      �                   p@���A��?J            �R@������������������������       �                     @�      �                   �v@
;&����?E            @Q@�      �                ��8�?؇���X�?             @������������������������       �                     @�      �                �:]�?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?V{q֛w�?>             O@�      �                PI�?�"U����?3            �I@�      �                   �?r�q��?             8@�      �                ����?      �?             (@������������������������       �                     @�      �                @��?���Q��?             @������������������������       �                      @�      �                   �@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                 �q�?�q�q�?             (@�      �                а2�?z�G�z�?
             $@�      �                   �?�����H�?	             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                ����?�<ݚ�?             ;@������������������������       �                      @�      �                ����?�����?             3@�      �                ����?      �?              @�      �                �8��?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                 /�?�C��2(�?             &@������������������������       �        	             "@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?���!pc�?             &@������������������������       �                     @�      �                   W�@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                ���?R�}e�.�?             :@�      �                �q�?R���Q�?             4@�      �                O�?�KM�]�?             3@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   ړ@�IєX�?             1@�      �                   �@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?�      �                   @�@�q�q�?             @������������������������       �                     @�      �                ��8�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   u�@4F�p�#�?�            �g@�      �                p�?$G$n��?%            �B@�      �                ��_�?��<b���?             7@�      �                ��8�?؇���X�?             5@�      �                   ��@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                   �?      �?             0@�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@������������������������       �                      @������������������������       �                     ,@�      �                   p�@:W��S��?�             c@�      �                p��?�	j*D�?4             J@�      �                ��8�? �o_��?2             I@�      �                ����?      �?             @������������������������       �                     �?������������������������       �                     @�      �                �V��?�5��
J�?.             G@������������������������       �                     �?�      �                   �@�<ݚ�?-            �F@������������������������       �                      @�      �                   �@����>�?%            �B@������������������������       �                     @�      �                  ���@H�V�e��?"             A@�      �                   �?�KM�]�?             3@�      �                 ���?����X�?             @�      �                   @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�      �                  �ɰ@�q�q�?             .@�      �                   �?      �?              @������������������������       �                     @�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�      �                 �	�?Fx$(�?d             Y@�      �                   �?�C��2(�?             &@������������������������       �        
             $@������������������������       �                     �?�                         4�@PN���?Y            @V@�             
             �?ȵHPS!�?             :@�      �                @��?z�G�z�?             .@�      �                   �?؇���X�?             ,@������������������������       �                     @�      �                P��?����X�?             @������������������������       �                     @�      �                @���?      �?             @������������������������       �                     �?�      �                   �?�q�q�?             @������������������������       �                     �?�      �                �q�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@                        �U�@p�EG/��??            �O@                      0���?      �?              @������������������������       �                     @������������������������       �                     �?      !                  �,�@��N`.�?7            �K@                       0��? �o_��?2             I@                        �̹@      �?0             H@	                         �?�����?&             C@
                      p��?�G��l��?             5@                        �*�@�	j*D�?             *@                        �|�@"pc�
�?             &@                      �Q>�?�����H�?	             "@������������������������       �                     @                      �q�?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         �?      �?              @������������������������       �                     @                         ?�@�q�q�?             @������������������������       �                     �?������������������������       �                      @                      ����?�t����?             1@������������������������       �                     �?                      ����?      �?             0@������������������������       �                     �?������������������������       �                     .@������������������������       �        
             $@������������������������       �                      @"      #                ��e�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @%      2                p���?������?             >@&      )                   �@d}h���?             <@'      (      
             �?      �?             @������������������������       �                     �?������������������������       �                     @*      1                �q�?      �?             8@+      0                   �?���}<S�?             7@,      -                � Q�?�q�q�?             @������������������������       �                     @.      /                �q�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@������������������������       �                     �?������������������������       �                      @4      �                �N�?�dG��?�           ؎@5      �                XUU�?������?@            �@6      �                �T�?�ՙ/�?�            `b@7      �                   �?�%�a�u�?�            �a@8      w                   �@ꟲ�4��?�            @a@9      f                   ��@�+Fi��?\             W@:      E                8\B ?�ɞ`s�?=            �N@;      >                    �@�����?             5@<      =                ��,?      �?              @������������������������       �                     �?������������������������       �                     �??      @                   �?�}�+r��?             3@������������������������       �                     *@A      B                ��d?r�q��?             @������������������������       �                     @C      D                   �?      �?              @������������������������       �                     �?������������������������       �                     �?F      Q                0��%?H�z�G�?(             D@G      H                    �@�q�q�?             .@������������������������       �                     @I      J                   (�@X�<ݚ�?	             "@������������������������       �                     @K      L                P�ԑ?�q�q�?             @������������������������       �                      @M      N                ��H#?      �?             @������������������������       �                     �?O      P                   u�@�q�q�?             @������������������������       �                      @������������������������       �                     �?R      S                   �? �o_��?             9@������������������������       �                     �?T      U                   @      �?             8@������������������������       �                     @V      W                   Pw@�q�q�?             2@������������������������       �                     �?X      ]                   �@�t����?             1@Y      \                   P�@      �?              @Z      [                   `�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @^      e                �E�?X�<ݚ�?	             "@_      d                   �?����X�?             @`      c                   �?�q�q�?             @a      b                    �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @g      l                P�ԑ?�P�*�?             ?@h      k                   �?8�Z$���?             *@i      j                  ��@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @m      t                   b�@b�2�tk�?             2@n      o                   @���Q��?
             $@������������������������       �                      @p      q                   �?      �?              @������������������������       �                     �?r      s                 ��?؇���X�?             @������������������������       �                     �?������������������������       �                     @u      v                   �?      �?              @������������������������       �                     @������������������������       �                     �?x      y                   �?��<b���?.             G@������������������������       �                     �?z      �                   �?z�G�z�?-            �F@{      �                  ��@ �Cc}�?             <@|      �                  ��@      �?             (@}      ~                   r�@"pc�
�?             &@������������������������       �                     @      �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@�      �                   ��@ҳ�wY;�?             1@������������������������       �                     @�      �                �W�'?��
ц��?             *@�      �                �|��?      �?              @�      �                   �?���Q��?             @������������������������       �                      @�      �                ��w?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                0�	�?��]��?�           h�@�      �                   g@�?�P�a�?,           �r@�      �                ����?X�<ݚ�?	             "@�      �                P��r?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                n��?��"��]�?#           0r@�      �                  �w�@ܷ��?��?"            r@�      �                ����?$C��_�?!           r@�      �                   �@bۘ�W^�?i            @Z@�      �                   A�@�9�a��?^            �W@�      �                   ��@����;�?]            @W@������������������������       �        	             "@�      �                   h�@��s����?T             U@������������������������       �                      @�      �                @`ރ?��r._�?R            �T@������������������������       �                     (@�      �                   l�@z�G�z�?F            �Q@�      �                ��8�?�r����?             >@�      �                   �?$�q-�?             :@������������������������       �                     2@�      �                0�	�?      �?              @������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @�      �                   զ@      �?(             D@������������������������       �                      @�      �                xǡ?���y4F�?&             C@������������������������       �                     �?�      �                @7�?��G���?%            �B@�      �                    �@      �?             @������������������������       �                      @������������������������       �                      @�      �                :�?6YE�t�?!            �@@�      �                   %�@��� ��?             ?@�      �                   �@      �?             (@�      �                �Po�?ףp=
�?
             $@������������������������       �                     �?������������������������       �        	             "@������������������������       �                      @�      �                   �?�}�+r��?             3@�      �                   �@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�      �                   �?���.�6�?�             g@�      �                PUU�?^�!~X�?5            �J@�      �                   �?��G���?%            �B@�      �                �jg�?      �?              @@�      �                   �?ףp=
�?             >@�      �                 ��?�nkK�?             7@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     4@�      �                   �?����X�?             @�      �                xǡ?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                 D)�?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                `~�?���Q��?             @�      �                ���?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     0@�      �                   �?؀���˲?�            ``@�      �                   ]�@�i�y�?~            �_@������������������������       �        2             I@�      �                   ��@�}�+r��?L             S@������������������������       �                     �?�      �                   ��@`2U0*��?K            �R@�      �                   ��@�����H�?             2@������������������������       �                     0@������������������������       �                      @�      �                   �?0�)AU��?9            �L@������������������������       �        0             H@�      �                ���?�����H�?	             "@�      �                ���?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                P�ԑ?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�                      �66�?4�2%ޑ�?�           x@�                      ����?|��?���?             ;@�                       ��}�?r�q��?             8@�      �                   �?�q�q�?             (@�      �                \��?�����H�?	             "@������������������������       �                     @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         p�@      �?             (@������������������������       �                      @                      ��
�?ףp=
�?
             $@������������������������       �                     @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @	      �                PUU�?,m�)6��?f           `v@
      g                   �?4��s?D�?J           �t@      T                ���?t�R2��?�            �k@      1                   �?fv�S��?�            �d@                      ��'�?R�(CW�?R            �T@                         �?�q�q�?             (@������������������������       �                     @                      Po�?�<ݚ�?	             "@                         �?      �?              @                         �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?      0                p��?(N:!���?F            �Q@                         �`@�θV�?E            @Q@������������������������       �                     �?      !      
             �?l��\��?D             Q@                         @��Y��]�?)            �D@������������������������       �                     >@                      ��.�?�C��2(�?             &@������������������������       �        	             "@                       `��?      �?              @������������������������       �                     �?������������������������       �                     �?"      /                   ��@�+$�jP�?             ;@#      ,                ��J�?�d�����?             3@$      +                   �?     ��?             0@%      &                   ԓ@�z�G��?
             $@������������������������       �                     @'      (                @��?և���X�?             @������������������������       �                      @)      *                   <�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @-      .                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?2      7                   �@��p �?R            �T@3      4                   @      �?              @������������������������       �                     @5      6                   �?      �?             @������������������������       �                     �?������������������������       �                     @8      Q                ��8�?����>�?J            �R@9      J                  ���@�q�q�?9            �L@:      C                   �?R���Q�?(             D@;      B                   �@ףp=
�?             >@<      A                   ��@      �?             (@=      >                p��?ףp=
�?
             $@������������������������       �                     @?      @                0*N�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     2@D      I                   �?���Q��?
             $@E      F                �?^�?�q�q�?             @������������������������       �                     @G      H                00��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @K      P                   й@j���� �?             1@L      O                 ���?����X�?             ,@M      N                   �@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @R      S                ����?�IєX�?             1@������������������������       �                     0@������������������������       �                     �?U      f                   �? ,��-�?;            �M@V      W                   ��@      �?              @@������������������������       �                     �?X      [                �^4�?��a�n`�?             ?@Y      Z                ����?      �?              @������������������������       �                     �?������������������������       �                     �?\      c                 �&�? 	��p�?             =@]      b                   �? 7���B�?             ;@^      a                   �?      �?              @_      `                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@d      e                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@h      i                ����?xZ�l ��?k            �Z@������������������������       �                      @j      �                   �?����X�?i            @Z@k      |                   �?>���Rp�?W            �U@l      w                �<t�?ZՏ�m|�?1            �H@m      t                   �?��(\���?(             D@n      o                   �?��?^�k�?#            �A@������������������������       �                     8@p      q                   �?�C��2(�?             &@������������������������       �                     @r      s                p��?      �?             @������������������������       �                     �?������������������������       �                     @u      v                @_r�?���Q��?             @������������������������       �                      @������������������������       �                     @x      {                  ���@X�<ݚ�?	             "@y      z                p}J�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @}      �                 ���?P����?&             C@~                      @��?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                p	��?���!pc�?!            �@@������������������������       �                     �?�      �                   �?      �?              @@�      �                   �@�t����?             1@������������������������       �                     �?�      �                ��k�?      �?             0@�      �                P{�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@�      �                �2�?���Q��?             .@�      �                   �?�q�q�?             @�      �                ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?�<ݚ�?	             "@������������������������       �                     �?�      �                �#��?      �?              @������������������������       �                     @�      �                ����?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                0���?      �?             2@������������������������       �                     @�      �                   �?X�Cc�?             ,@������������������������       �                     @�      �                �k��?X�<ݚ�?	             "@�      �                ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     <@�      �                ��J�?b�MKm�?�            `c@�      �                �rv�?����5�?=            �N@�      �                   �?�E��ӭ�?6             K@�      �                   �@��S���?             .@�      �                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�      �                 ��?      �?              @������������������������       �                     �?������������������������       �                     @�      �                ���?:�&���?'            �C@�      �                ��?ҳ�wY;�?             1@�      �                �8��?������?             .@������������������������       �                     @�      �                @��?      �?              @������������������������       �                      @�      �                І��?�q�q�?             @������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                   �?���7�?             6@������������������������       �                     .@�      �                PUU�?؇���X�?             @�      �                ��8�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                �8��?����X�?             @������������������������       �                      @������������������������       �                     @�      �                 R��?@�҇��?^            �W@�      �                �ۋ�?���*~�?Y            @V@�      �                �q�?����X�?8             L@�      �                0=P�?�q�q��?0             H@�      �                   �?��S�ۿ?             .@������������������������       �                     &@�      �                0)��?      �?             @������������������������       �                     �?������������������������       �                     @�      �                ���?:ɨ��?!            �@@�      �                �q�?և���X�?             5@�      �                   @�t����?             1@�      �                   �?      �?             0@�      �                  ���@���Q��?
             $@�      �                   ��@      �?              @������������������������       �                     �?�      �                �8��?؇���X�?             @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?�8��8��?             (@������������������������       �        	             "@�      �      
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                P��?      �?              @������������������������       �                     @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   �@�C��2(�?!            �@@�      �                p��?      �?              @@������������������������       �                     1@�      �                   �?�r����?             .@�      �                   �?      �?              @�      �                   �?؇���X�?             @�      �                Pu��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                P�?�M���?�	           �@�      �                   �?،(��?�           �@�      \                   �?x��ėb�?w           ��@�      1                �ae�?P;ߣ	H�?|           ��@�                        �Fa? �t��̮?�           0|@�      �                �J_?z�G�z�?
             $@�      �                   �?�����H�?	             "@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?            	             �?P����?�           �{@                      ����?�U�=���?B            �P@������������������������       �                     �?                        ���@����?A            @P@                         8�@�����?*             E@                         �?��p\�?)            �D@                         �?�}�+r��?&             C@������������������������       �                     8@	      
                   �?؇���X�?             ,@������������������������       �        	             "@                         �?���Q��?             @������������������������       �                      @������������������������       �                     @                      ��/�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     7@                         8x@�v¢?w           pw@                         t@؇���X�?             ,@                         �?$�q-�?             *@������������������������       �                     &@                       oc�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                       �8��?�A����?i           �v@                      �Fj�?�J�Է�?�            �n@                      �X�?`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?������������������������       �        �            `k@!      "                   �?ȑ����?u            @]@������������������������       �                     �?#      0                   �? �^�@̩?t             ]@$      /                p;{�?����˵�?;            �M@%      .                 �a�?l��\��?"             A@&      '                �ئ�?�FVQ&�?!            �@@������������������������       �                     1@(      )                �yj�?      �?             0@������������������������       �                     �?*      +                PUU�?��S�ۿ?             .@������������������������       �                     &@,      -                @��?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     9@������������������������       �        9            �L@2      ;                ���?�L���?�             g@3      :                ���?�	j*D�?             *@4      5                p�Ǽ?"pc�
�?             &@������������������������       �                     �?6      7                   �?ףp=
�?
             $@������������������������       �                      @8      9                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @<      Q                �8��?�Ts�k��?�            �e@=      P                Ё��?t�U����?C            �P@>      A                   �@��IF�E�?B            �P@?      @                   �m@      �?             @������������������������       �                      @������������������������       �                      @B      M                ����?6uH���?>             O@C      H                   @�h����?8             L@D      E                �[�?����?�?-            �F@������������������������       �        '            �C@F      G                0j��?r�q��?             @������������������������       �                     �?������������������������       �                     @I      J                   �?"pc�
�?             &@������������������������       �                     @K      L                ��8�?      �?             @������������������������       �                      @������������������������       �                      @N      O                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?R      S                �$��?��?^�k�?i            @Z@������������������������       �        V            �U@T      U                   �?�S����?             3@������������������������       �                     (@V      W                ��E�?և���X�?             @������������������������       �                      @X      [                09y�?z�G�z�?             @Y      Z                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @]      f                �	��?�vps�?�            `o@^      a                   �@�q�q�?             5@_      `                ��S�?r�q��?             @������������������������       �                     �?������������������������       �                     @b      c                   �?�r����?             .@������������������������       �                     �?d      e                   ٸ@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?g      h                    8@���AY5�?�            �l@������������������������       �                     �?i      r                �t:�?�p5]y�?�            �l@j      k                �0@�?�g�y��?>             O@������������������������       �        6             K@l      m                �o�?      �?              @������������������������       �                     �?n      o                   �?؇���X�?             @������������������������       �                     @p      q                   گ@      �?              @������������������������       �                     �?������������������������       �                     �?s      v                �̱�?~n��W��?�            �d@t      u                0��?      �?             @������������������������       �                     �?������������������������       �                     @w      �                  �u�@�Ǐ�?�            `d@x      {                �q�?K�|%��?}            @_@y      z                �D�?�q�q�?             @������������������������       �                      @������������������������       �                     �?|      �                  �´@��.��?z            �^@}      �                pff�?�io�?t             ]@~      �                pt3�?0�W���?e            @Y@      �                   �R@�J�4�?d             Y@������������������������       �                     �?�      �                ����?6YE�t�?c            �X@�      �                Ц��?�r����?Z            �V@�      �                p+��?�3Ea�$�?.             G@�      �      
             �?��a�n`�?             ?@������������������������       �                     2@�      �                   �?�θ�?             *@������������������������       �                     @�      �                   c�@և���X�?             @������������������������       �                     @�      �      	             �?      �?             @������������������������       �                     @������������������������       �                     �?�      �                �_=�?���Q��?             .@������������������������       �                      @�      �                   �?�	j*D�?             *@�      �                ����?X�<ݚ�?	             "@�      �                   �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                p��?t��ճC�?,             F@������������������������       �                     5@�      �                p�#�?�LQ�1	�?             7@�      �                   ��@�C��2(�?             6@������������������������       �                     �?�      �                �8��?���N8�?             5@�      �                   ��@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@������������������������       �                     �?�      �                0���?�q�q�?	             "@�      �                   �@���Q��?             @�      �                �q�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�      �      	             �?      �?             @������������������������       �                     @������������������������       �                     @�      �                  ���@P�Lt�<�?&             C@������������������������       �                     <@�      �                  �ʹ@ףp=
�?
             $@������������������������       �                     �?������������������������       �        	             "@�      �                0���? @ެ[�?           @�@�      �                ���? D�R��?3           ��@�      �                PHy�?����3�?1           ��@�      �                �q�?�����?�            �@�      �                PUU�?��Vl��?�           `{@�      �                  � �@�:!�g��?X           �u@������������������������       �        �            �o@�      �                   *�@hl �&�?\             W@������������������������       �                     �?�      �                   �?p�C��?[            �V@������������������������       �        A            @P@�      �                �(�?$�q-�?             :@�      �                ���?      �?              @�      �                   �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�      �                   h�@`�q�0ܴ?^            �W@�      �                   ܅@8�Z$���?             *@�      �                0��?�8��8��?             (@�      �                ��׽?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             $@������������������������       �                     �?�      �                @��?F|/ߨ�?Q            @T@�      �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?�"w����?L             S@�      �                ���?�����H�?	             "@������������������������       �                     �?������������������������       �                      @������������������������       �        C            �P@�      �      	             �? ��e{?*           �r@�      �                p��?XB���?             =@������������������������       �                     ;@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                   �p@�      �                 ��? 7���B�?Q            @T@������������������������       �                     �?�      �      
             �?�(\����?P             T@�      �                �"X�?�t����?             1@������������������������       �                     �?�      �                   �?      �?             0@�      �                `UU�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �        ?            �O@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        �            �k@�      ~                   �?r�q��?p           ��@�      y                �N�?�+e�X�?E           Pt@�      x                PUU�?�t����??           �s@�                      ���?Z�/�j��?*           �r@�                         ��@������?[            �V@�                          �@�+e�X�?2             I@�                      �q�?���c�H�?1            �H@�      �                @��?�3Ea�$�?.             G@�      �                @���?���Q��?
             $@������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                   @4?,R��?$             B@�      �                    �@���7�?             6@�      �                   �z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�            	             �?����X�?             ,@�                      �k��?և���X�?             @                          �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?	                      P�c�?��p\�?)            �D@
                      p"=�?�<ݚ�?	             "@������������������������       �                     @                      Cw�?�q�q�?             @������������������������       �                     �?������������������������       �                      @                      �7��?      �?              @@                        �<�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@      ]                `q'�?�m淣�?�            �i@      >                p��?�X���?�            �`@      %                   �?���mC�?U            @U@      $                   �?r�q��?             8@      !                mQ�?�G�z��?             4@                       ��?�n_Y�K�?             *@������������������������       �                      @                         Q�@���!pc�?             &@������������������������       �                      @                       ���?�����H�?	             "@                      ��8�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @"      #                   ��@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @&      '                p��?`��:�?=            �N@������������������������       �                     ,@(      )                   �}@�*/�8V�?/            �G@������������������������       �                      @*      3      
             �?�<ݚ�?-            �F@+      ,                @��?b�2�tk�?             2@������������������������       �                     @-      .                   :�@d}h���?             ,@������������������������       �                      @/      0                p���?      �?             @������������������������       �                      @1      2                   �?      �?             @������������������������       �                     @������������������������       �                     �?4      ;                   �@�����H�?             ;@5      6                   �?HP�s��?             9@������������������������       �                     0@7      :                0���?�<ݚ�?	             "@8      9                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @<      =                ��8�?      �?              @������������������������       �                     �?������������������������       �                     �??      N      	             �?JJ����?/            �G@@      E                   �?�û��|�?             7@A      B                ����?�����H�?	             "@������������������������       �                     @C      D                   �?      �?              @������������������������       �                     �?������������������������       �                     �?F      G                   �?և���X�?             ,@������������������������       �                     @H      I                ����?���Q��?
             $@������������������������       �                     @J      M                ��k�?և���X�?             @K      L                ���?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @O      \                ����?�q�q�?             8@P      Q                 ���?���!pc�?             6@������������������������       �                     @R      S                Pc�?      �?             0@������������������������       �                     @T      U                   `\@�θ�?             *@������������������������       �                     �?V      W                `UU�?r�q��?             (@������������������������       �                     @X      [                 �1�?�q�q�?             @Y      Z                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @^      q                `4O�?��n�?K            �R@_      p      	             �?؇���X�??            �O@`      a                   �@�θ�?'            �C@������������������������       �        	             "@b      e                   m�@�z�G��?             >@c      d                ���?      �?             @������������������������       �                     �?������������������������       �                     @f      g                  �հ@�θ�?             :@������������������������       �        	             "@h      i                   ۱@ҳ�wY;�?             1@������������������������       �                     @j      m                   �?d}h���?             ,@k      l                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @n      o                �q�?�C��2(�?             &@������������������������       �        
             $@������������������������       �                     �?������������������������       �                     8@r      s                Pq��?�q�q�?             (@������������������������       �                     @t      w                ����?      �?              @u      v      
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     5@z      }                   �?�q�q�?             @{      |                0�N�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @      �                ��,�?���}<S�?+           �r@�      �                p۶�?���Q��?             @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                p��?��v�u�?&           `r@�      �                `���?pb����?�             g@�      �                 �J�?p�qG�?`             X@�      �                   B�@r�q��?             8@�      �                ���?�LQ�1	�?             7@�      �                �rv�?�C��2(�?             6@�      �                ����?���N8�?             5@������������������������       �                     1@�      �                ��~�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                �_��?�k~X��?H             R@�      �                 �p�?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �        9            �L@�      �                p�#�?NKF����?Y            @V@�      �                �8��?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                ��8�?0,Tg��?T             U@�      �                0��?����X�?             <@�      �                   �?"pc�
�?             6@������������������������       �        	             "@�      �                0���?�	j*D�?             *@�      �                ��`�?      �?              @������������������������       �                      @�      �                 5�?�q�q�?             @������������������������       �                     �?�      �                 ��?z�G�z�?             @������������������������       �                     @�      �                �1�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                   �?4և����?8             L@�      �                 .�?     ��?             0@�      �                p��?�r����?             .@�      �                p���?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             $@������������������������       �                     �?�      �                   ��@P���Q�?(             D@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                0���?�?�|�?%            �B@������������������������       �                     ;@�      �                `���?ףp=
�?
             $@������������������������       �                     �?������������������������       �        	             "@�      �                 �>�?��wڝ�?m            @[@�      �                P�?�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?������������������������       �        Z            �V@��|      �t�b�values�hhK ��h��R�(KM�KK��hu�B0|       *�@     `�@     ��@     ��@      �@     ��@      w@     �@     �i@      i@      c@      g@     �O@     �Z@     �H@     �P@     �H@      M@     �G@     �G@      D@      G@     �A@     �F@      9@      7@      8@      0@      .@      @      �?       @      �?                       @      ,@       @       @       @      @              @       @      �?       @      �?                       @       @              @              "@      (@       @              @      (@      �?      @              @      �?       @               @      �?              @      @      @              @      @       @      @       @      �?       @                      �?              @      �?              �?      @              @      �?              $@      6@      @      5@      @      3@       @      3@              (@       @      @      �?              �?      @      �?      �?              �?      �?                      @      �?              @       @      �?       @      �?                       @       @              @      �?      @                      �?      @      �?              �?      @              @      �?      @                      �?       @      &@       @      @      �?      @              @      �?       @      �?                       @      �?                      @               @      ,@      D@      @      A@      �?              @      A@      @      A@      @      ?@              5@      @      $@      �?      $@               @      �?       @               @      �?               @               @      @               @       @      �?       @                      �?      �?              @      @      @              @      @      �?      @              @      �?      �?              �?      �?               @             �V@     �S@     �V@      R@     �T@     �M@     �D@     �C@      >@      B@      2@      $@      *@      @      *@       @      *@      �?      *@                      �?              �?              �?      @      @      @      @      �?      @              @      �?               @               @              (@      :@              @      (@      5@       @              $@      5@       @      &@      @      &@      @      @      @      @      @       @               @      @                      @       @                      @      @               @      $@              $@       @              &@      @               @      &@      �?      "@               @      �?              �?       @              E@      4@      8@      @              �?      8@      @       @              0@      @      0@      @       @      @       @       @       @      �?       @                      �?              �?               @       @                      �?      2@      ,@              @      2@      "@      1@      @      .@       @      .@      �?       @      �?              �?       @              *@                      �?       @      @       @      �?       @                      �?               @      �?      @              @      �?              @      *@      @      �?      @                      �?       @      (@      �?      (@      �?                      (@      �?                      @     �J@      0@      J@      &@      <@      $@      1@      $@      1@      @      &@      �?      $@              �?      �?              �?      �?              @      @       @      @      �?              �?      @              @      �?      �?      �?                      �?      @      �?      �?      �?              �?      �?              @                      @      &@              8@      �?      4@              @      �?      @                      �?      �?      @      �?                      @     �d@     �{@      9@     �b@              ?@      9@      ^@      .@     �C@      @      ?@      �?              @      ?@      �?              @      ?@              *@      @      2@      �?              @      2@      �?      �?      �?                      �?       @      1@              (@       @      @       @      �?       @                      �?              @      "@       @       @      @              �?       @      @       @       @      @       @      �?       @      �?                       @       @              @                      �?      �?      @              @      �?              $@     @T@      @      2@              $@      @       @      @       @       @       @              @       @      �?              �?       @               @               @              @     �O@      �?     �B@              @@      �?      @      �?                      @      @      :@      �?               @      :@       @      *@      �?      *@      �?      @              @      �?                      "@      �?                      *@     `a@      r@     �O@     �Q@     �C@     �K@      @      1@       @      .@      �?      ,@              $@      �?      @              @      �?      �?      �?                      �?      �?      �?      �?                      �?      @       @      �?       @               @      �?               @              A@      C@      ?@      C@      ?@      @@      8@      3@      @              2@      3@       @      ,@              @       @      @               @       @      @      @              @      @              @      @       @               @      @              $@      @      @      �?       @      �?       @                      �?      @              @      @      @      �?              �?      @                      @      @      *@      @      *@      @      *@      @      @              @      @      @      @              �?      @              @      �?                      @      �?               @                      @      @              8@      0@      $@      *@      @              @      *@      @      @      @      @              @      @      �?      @                      �?       @              �?       @      �?       @      �?                       @              @      ,@      @      ,@       @      (@               @       @       @                       @              �?      S@     `k@     �G@     �W@       @      9@      �?      7@      �?      @              @      �?                      1@      �?       @      �?                       @     �F@     �Q@      "@       @               @      "@              B@      Q@     �A@     �L@      >@      L@      *@      B@      $@      *@      @      $@      �?      "@               @      �?      �?              �?      �?               @      �?       @                      �?      @      @      @              �?      @              @      �?              @      7@              3@      @      @      @      �?      @                      �?              @      1@      4@      @              (@      4@      �?      "@      �?      �?      �?                      �?               @      &@      &@              @      &@       @      @       @               @      @              @      @       @      @              @       @               @              @      �?      @                      �?      �?      &@              &@      �?              =@      _@      @              :@      _@      8@     �^@      7@     �^@      2@     �\@      *@     �K@      "@      4@       @      (@      @      (@      @      @      @       @      @                       @               @               @      @              �?       @      �?       @               @      �?                      @      @     �A@       @      @       @      �?              �?       @                      @       @      >@      �?      <@              6@      �?      @              @      �?              �?       @               @      �?              @     �M@              9@      @      A@      �?              @      A@              2@      @      0@       @      �?       @                      �?       @      .@      �?      �?              �?      �?              �?      ,@      �?      @              @      �?                      &@      @      "@      @      "@      �?               @      "@              @       @       @      �?              �?       @      �?                       @       @              �?               @      �?       @                      �?     p�@     �z@     `k@     �M@     �S@     �A@               @     �S@     �@@      8@      @      @      @       @      @       @      �?              �?       @                       @      @              1@             �K@      >@      B@      ;@      7@      $@      @      @      @       @      @              �?       @               @      �?              �?      @              @      �?              1@      @      ,@      �?              �?      ,@              @       @               @      @              *@      1@              @      *@      (@      @      "@      @      "@              @      @      @               @      @      �?      @                      �?       @               @      @      @               @      @              @       @              3@      @              �?      3@       @      .@              @       @      @              �?       @               @      �?             �a@      8@      J@      1@      ?@      @       @      @               @       @      �?       @                      �?      =@       @      2@              &@       @              �?      &@      �?      �?      �?      �?                      �?      $@              5@      (@      2@      @      &@      @      "@      �?       @              �?      �?      �?                      �?       @      @      �?              �?      @              @      �?              @              @      @      @                      @      V@      @      O@       @     �G@              .@       @      ,@              �?       @               @      �?              :@      @      :@      @      $@              0@      @      @      @       @              �?      @              @      �?              *@      �?      �?      �?              �?      �?              (@                      �?     0{@     0w@     �g@     �[@      c@     @R@     �W@     �N@     �J@     �H@     �H@     �A@     �A@     �@@     �@@      5@      @      @      @                      @      >@      ,@      ,@      *@      @      �?      @               @      �?       @                      �?      @      (@      @      @      �?      @              @      �?              @      �?      @                      �?              @      0@      �?       @      �?              �?       @              ,@               @      (@      �?              �?      (@      �?      �?              �?      �?                      &@      ,@       @      &@              @       @      @                       @      @      ,@              *@      @      �?              �?      @             �D@      (@      @      @              @      @      �?      @                      �?     �B@       @      @@      @       @      @       @      �?              �?       @                       @      8@      �?      @      �?      @                      �?      5@              @      @      @      �?              �?      @                      @     �M@      (@     �F@      @      7@      @      6@      @      *@              "@      @              �?      "@       @              �?      "@      �?      @               @      �?              �?       @              �?       @               @      �?              6@      �?      @      �?      @                      �?      0@              ,@      @      @      @      �?      @              @      �?              @      �?      @                      �?      "@      �?      �?      �?      �?                      �?       @             �A@      C@      .@       @      @      @              @      @       @      �?       @      �?                       @       @              (@      @      @      @      @              �?      @              @      �?              @              4@      >@       @      $@      �?              �?      $@              "@      �?      �?      �?                      �?      2@      4@      @              *@      4@              @      *@      ,@      "@      @      �?      @              @      �?               @      �?      @              �?      �?              �?      �?              @      $@      �?      "@      �?                      "@      @      �?      @                      �?     �n@     @p@      L@      <@      =@       @      *@      @               @      *@      @      @              @      @      �?      @      �?                      @      @      �?      �?      �?      �?                      �?      @              0@      �?              �?      0@              ;@      4@      0@       @      ,@      @      ,@      @      (@      �?      �?      �?              �?      �?              &@               @       @       @                       @              �?       @      @              @       @      �?       @                      �?      &@      (@              @      &@      "@      @              @      "@       @      @              @       @       @       @                       @      @      @      @              �?      @      �?                      @     �g@      m@      <@     �P@      ,@      $@              @      ,@      @      @              "@      @               @      "@      @       @       @      @               @       @               @       @              �?      @              @      �?              ,@      L@      �?      =@      �?      @              @      �?                      9@      *@      ;@      @              $@      ;@      "@      ,@       @      "@      �?              �?      "@      �?      �?      �?                      �?               @      @      @      @      �?      �?      �?      �?                      �?      @              �?      @              @      �?              �?      *@              &@      �?       @               @      �?             `d@     �d@     �a@     �c@      O@      H@     �L@      H@      C@     �D@      @             �@@     �D@              @     �@@      B@      @      �?      @              �?      �?      �?                      �?      ;@     �A@      3@      @@      *@      &@      "@      @      @               @      @               @       @      �?              �?       @              @       @       @       @      �?       @               @      �?              �?               @              @      5@               @      @      *@      @      @      @      �?              �?      @                       @      �?      $@              "@      �?      �?              �?      �?               @      @      @               @      @              @       @              3@      @      1@      @      1@       @      �?      �?              �?      �?              0@      �?      @      �?      @                      �?      (@                      �?       @      @              @       @      �?              �?       @              @             �S@     �[@      @      @@      @      2@      @      2@       @      @              @       @              �?      .@      �?      @              @      �?                      (@       @                      ,@     �R@     �S@      B@      0@      B@      ,@      �?      @      �?                      @     �A@      &@              �?     �A@      $@       @              ;@      $@              @      ;@      @      1@       @      @       @      @      �?      @                      �?              �?      (@              $@      @      @      @              @      @      �?              �?      @              @                       @      C@      O@      $@      �?      $@                      �?      <@     �N@      @      7@      @      (@       @      (@              @       @      @              @       @       @      �?              �?       @              �?      �?      �?      �?                      �?      �?                      &@      9@      C@      @      �?      @                      �?      2@     �B@      ,@      B@      (@      B@      (@      :@      $@      &@      @      "@       @      "@      �?       @              @      �?       @      �?                       @      �?      �?      �?                      �?       @              @       @      @              �?       @      �?                       @       @      .@      �?              �?      .@      �?                      .@              $@       @              @      �?              �?      @              6@       @      6@      @      �?      @      �?                      @      5@      @      5@       @      @       @      @              �?       @      �?                       @      1@                      �?               @     @�@     `n@     h�@     `f@     �V@      L@     �V@     �I@     �V@     �G@     �K@     �B@      E@      3@      3@       @      �?      �?              �?      �?              2@      �?      *@              @      �?      @              �?      �?      �?                      �?      7@      1@      @      $@              @      @      @      @               @      @               @       @       @      �?              �?       @               @      �?              2@      @              �?      2@      @      @              (@      @              �?      (@      @      @      �?      @      �?      @                      �?      @              @      @      @       @      �?       @      �?      �?              �?      �?                      �?      @                       @      *@      2@       @      &@       @      @              @       @                       @      &@      @      @      @       @               @      @      �?              �?      @      �?                      @      @      �?      @                      �?      B@      $@              �?      B@      "@      9@      @      "@      @      "@       @      @              @       @               @      @                      �?      0@              &@      @      @              @      @      @      @      @       @       @              �?       @               @      �?                      @      @      �?              �?      @                      @              @     ��@     �^@     �p@     �A@      @      @       @      @       @                      @      @             @p@      ?@     @p@      >@     @p@      =@      V@      1@     @S@      1@     @S@      0@      "@              Q@      0@               @      Q@      ,@      (@              L@      ,@      :@      @      8@       @      2@              @       @      @              �?       @      �?                       @       @       @               @       @              >@      $@               @      >@       @              �?      >@      @       @       @               @       @              <@      @      ;@      @      "@      @      "@      �?              �?      "@                       @      2@      �?      @      �?      @                      �?      .@              �?      �?              �?      �?                      �?      &@             �e@      (@      G@      @      >@      @      <@      @      ;@      @      6@      �?       @      �?              �?       @              4@              @       @      �?       @      �?                       @      @              �?      �?              �?      �?               @      @       @      �?              �?       @                       @      0@             �_@      @     �^@      @      I@              R@      @              �?      R@      @      0@       @      0@                       @      L@      �?      H@               @      �?      �?      �?      �?                      �?      @              @      �?              �?      @                      �?              �?     �r@      V@      *@      ,@      *@      &@      @       @      �?       @              @      �?      �?              �?      �?              @              "@      @               @      "@      �?      @               @      �?              �?       @                      @     �q@     �R@      p@     �R@     �f@      E@     �_@      C@     @Q@      *@      @      @              @      @       @      @      �?      �?      �?      �?                      �?      @                      �?      O@       @      O@      @              �?      O@      @      D@      �?      >@              $@      �?      "@              �?      �?              �?      �?              6@      @      ,@      @      *@      @      @      @      @              @      @               @      @      �?              �?      @              @              �?       @      �?                       @       @                      �?     �L@      9@      @      @              @      @      �?              �?      @              K@      4@      C@      3@      ?@      "@      ;@      @      "@      @      "@      �?      @              @      �?              �?      @                       @      2@              @      @      @       @      @              �?       @               @      �?                      @      @      $@      @      $@      @      @      @                      @              @      @              0@      �?      0@                      �?     �K@      @      <@      @              �?      <@      @      �?      �?      �?                      �?      ;@       @      :@      �?      @      �?      @      �?      @                      �?      @              3@              �?      �?              �?      �?              ;@             �R@      @@               @     �R@      >@     �P@      5@     �D@       @     �B@      @      A@      �?      8@              $@      �?      @              @      �?              �?      @              @       @               @      @              @      @      @      �?              �?      @                      @      9@      *@      �?      @              @      �?              8@      "@              �?      8@       @      .@       @              �?      .@      �?       @      �?       @                      �?      *@              "@      @       @      @      �?      @      �?                      @      �?              @       @              �?      @      �?      @              �?      �?      �?                      �?      "@      "@              @      "@      @      @              @      @      @      �?              �?      @                      @      <@             �V@      P@      4@     �D@      .@     �C@       @      @      �?      @      �?                      @      @      �?              �?      @              @      @@      @      &@      @      &@              @      @      @       @               @      @              @       @      �?       @                      �?       @              �?      5@              .@      �?      @      �?      �?              �?      �?                      @      @       @               @      @             �Q@      7@     �Q@      3@      D@      0@     �B@      &@      ,@      �?      &@              @      �?              �?      @              7@      $@      (@      "@      (@      @      (@      @      @      @      @       @              �?      @      �?      @              �?      �?      �?                      �?               @      @                      �?              @      &@      �?      "@               @      �?              �?       @              @      @              @      @      �?      @                      �?      >@      @      >@       @      1@              *@       @      @       @      @      �?       @      �?       @                      �?      @                      �?      @                      �?      �?      @              @      �?             ��@     �f@     �@     @S@     ��@     @P@     ��@      =@     P{@      ,@       @       @       @      �?      �?      �?              �?      �?              @                      �?     �z@      (@     �N@      @              �?     �N@      @      C@      @      C@      @      B@       @      8@              (@       @      "@              @       @               @      @               @      �?              �?       @                      �?      7@              w@      @      (@       @      (@      �?      &@              �?      �?      �?                      �?              �?     @v@      @     `n@      �?      8@      �?      8@                      �?     `k@             @\@      @              �?     @\@      @      L@      @      ?@      @      ?@       @      1@              ,@       @              �?      ,@      �?      &@              @      �?              �?      @                      �?      9@             �L@             @e@      .@      "@      @      "@       @              �?      "@      �?       @              �?      �?              �?      �?                       @      d@      &@     �M@       @     �M@      @       @       @       @                       @     �L@      @     �J@      @      F@      �?     �C@              @      �?              �?      @              "@       @      @               @       @               @       @              @       @      @                       @              �?     �Y@      @     �U@              0@      @      (@              @      @               @      @      �?      �?      �?      �?                      �?      @             �j@      B@      ,@      @      �?      @      �?                      @      *@       @              �?      *@      �?      *@                      �?      i@      =@              �?      i@      <@      N@       @      K@              @       @              �?      @      �?      @              �?      �?      �?                      �?     �a@      :@      �?      @      �?                      @     �a@      7@     �Y@      6@      �?       @               @      �?             �Y@      4@     �X@      1@      U@      1@      U@      0@              �?      U@      .@     �S@      (@     �B@      "@      <@      @      2@              $@      @      @              @      @      @              �?      @              @      �?              "@      @               @      "@      @      @      @      @      �?      @                      �?              @      @             �D@      @      5@              4@      @      4@       @              �?      4@      �?      @      �?              �?      @              0@                      �?      @      @       @      @       @      �?       @                      �?               @      @                      �?      .@              @      @              @      @             �B@      �?      <@              "@      �?              �?      "@             �@      (@     8�@      (@     0�@      &@     ��@       @     �z@      @     Pu@      @     �o@             @V@      @              �?     @V@       @     @P@              8@       @      @       @      �?       @               @      �?              @              2@             �V@      @      &@       @      &@      �?      �?      �?      �?                      �?      $@                      �?     �S@       @      @      �?      @                      �?     �R@      �?       @      �?              �?       @             �P@             �r@      �?      <@      �?      ;@              �?      �?              �?      �?             �p@             �S@      @              �?     �S@       @      .@       @              �?      .@      �?       @      �?              �?       @              *@             �O@              �?      �?              �?      �?             �k@             @�@      Z@     �n@     �S@     �n@     �R@      l@     �R@      S@      .@      C@      (@      C@      &@     �B@      "@      @      @      @               @      @              @       @              ?@      @      5@      �?      @      �?      @                      �?      2@              $@      @      @      @      @      �?              �?      @                      @      @              �?       @               @      �?                      �?      C@      @      @       @      @              �?       @      �?                       @      ?@      �?      �?      �?      �?                      �?      >@             �b@     �M@     �U@     �F@      O@      7@      *@      &@      "@      &@       @      @               @       @      @               @       @      �?      �?      �?      �?                      �?      @              �?      @      �?                      @      @             �H@      (@      ,@             �A@      (@               @     �A@      $@      &@      @              @      &@      @       @              @      @       @              �?      @              @      �?              8@      @      7@       @      0@              @       @      �?       @      �?                       @      @              �?      �?      �?                      �?      9@      6@      "@      ,@      �?       @              @      �?      �?      �?                      �?       @      @      @              @      @              @      @      @      @      �?              �?      @                       @      0@       @      0@      @      @              $@      @              @      $@      @              �?      $@       @      @              @       @      �?       @      �?                       @      @                       @     �N@      ,@      K@      "@      >@      "@      "@              5@      "@      �?      @      �?                      @      4@      @      "@              &@      @              @      &@      @      �?       @      �?                       @      $@      �?      $@                      �?      8@              @      @      @              @      @      �?      @      �?                      @       @              5@               @      @       @      �?       @                      �?              @     q@      :@       @      @       @      �?       @                      �?               @     �p@      7@     `d@      6@     �V@      @      4@      @      4@      @      4@       @      4@      �?      1@              @      �?              �?      @                      �?              �?              �?     �Q@      �?      ,@      �?      ,@                      �?     �L@              R@      1@      �?      @      �?                      @     �Q@      *@      4@       @      2@      @      "@              "@      @      @      @       @               @      @      �?              �?      @              @      �?      �?      �?                      �?      @               @      @              @       @             �I@      @      *@      @      *@       @      @       @      @                       @      $@                      �?      C@       @       @      �?              �?       @              B@      �?      ;@              "@      �?              �?      "@              [@      �?      2@      �?      2@                      �?     �V@        �t�bub�_sklearn_version��1.2.2�ub.