��5      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�K*�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�gender��SeniorCitizen��Partner��
Dependents��tenure��PhoneService��MultipleLines��InternetService��OnlineSecurity��OnlineBackup��DeviceProtection��TechSupport��StreamingTV��StreamingMovies��Contract��PaperlessBilling��PaymentMethod��MonthlyCharges��TotalCharges�et�b�n_features_in_�K�
n_outputs_�K�classes_�hhK ��h��R�(KK��h �i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�h�scalar���hDC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��hD�C       �t�bK��R�}�(h	K�
node_count�M��nodes�hhK ��h��R�(KM���h �V56�����R�(Kh$N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hfh �i8�����R�(KhENNNJ����J����K t�bK ��hghqK��hhhqK��hih �f8�����R�(KhENNNJ����J����K t�bK��hjhxK ��hkhqK(��hlhxK0��uK8KKt�b�B��        �                   �?���%���?           �@       �                   �?n��"O�?           �@       l                ����?H6�(���?0           `�@                          �?~��6��?�           ��@       �                 �|�?XK�~���?�           py@                        �Ӻ}?�j4����?R            u@       ^                 �Ӻm?l��@���?�             e@       ]                    �?��|��L�?s            �\@	       T                    �?���
��?k            �Z@
       O                    �?      �?^            �W@       L       	             �?v ��?V            �U@       5                 `��?     ��?P             T@       2                    �?�q���?0             H@                           �?���Q��?(             D@                        �09h?      �?             4@                        0�h?     ��?             0@                         ��G?d}h���?             ,@                           @���Q��?             @������������������������       �                      @������������������������       �                     @                           @�����H�?	             "@������������������������       �                     @                        XUU�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @       )                   �?�G�z��?             4@       (                 �dı?�z�G��?
             $@       '                    �?և���X�?             @                         0&�D?�q�q�?             @������������������������       �                     �?!       "                 ��DE?���Q��?             @������������������������       �                     �?#       &                     �?      �?             @$       %                 ���G?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @*       -                     �?���Q��?
             $@+       ,                 �
n�?      �?             @������������������������       �                     �?������������������������       �                     @.       1                 ��h?r�q��?             @/       0                 ���g?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @3       4                    �?      �?              @������������������������       �                     @������������������������       �                     �?6       I                    �?     ��?              @@7       B                 @5�?�<ݚ�?             ;@8       9                    @��2(&�?             6@������������������������       �                     &@:       A                 ���i?���!pc�?             &@;       @                  /��?և���X�?             @<       ?                    �?�q�q�?             @=       >                 0��h?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @C       H                     �?���Q��?             @D       E                 �`�m?�q�q�?             @������������������������       �                     �?F       G                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @J       K                 �^!�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @M       N                 82��?r�q��?             @������������������������       �                     �?������������������������       �                     @P       Q                 p���?      �?              @������������������������       �                     @R       S                    @      �?              @������������������������       �                     �?������������������������       �                     �?U       \                  �ih?8�Z$���?             *@V       [                 p@��?      �?              @W       X       	             �?؇���X�?             @������������������������       �                     @Y       Z                  �8U?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @_       v                 @؋�?������?6             K@`       e                 ��p?��r._�?)            �D@a       b                    �?      �?             0@������������������������       �                     *@c       d                 ���?�q�q�?             @������������������������       �                      @������������������������       �                     �?f       s       	             �?�+e�X�?             9@g       l                 �� �?"pc�
�?             6@h       k                  ʣ�?�8��8��?             (@i       j                 ��y?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             "@m       n                 P�n�?�z�G��?
             $@������������������������       �                      @o       r                 ���p?      �?              @p       q       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @t       u                  C��?�q�q�?             @������������������������       �                     �?������������������������       �                      @w       x                  ��?��
ц��?             *@������������������������       �                     @y       ~                  ��t?�q�q�?	             "@z       {                    �?؇���X�?             @������������������������       �                     @|       }                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                 ��8�?|ƀQK��?�             e@�       �       
             �?X�<ݚ�?�            @d@�       �                 @؋�?���A��?�            �a@�       �                 @���?vs�G��?v            �]@�       �                    �?r�z-��?5            �J@�       �                 ����?�q�q�?             8@�       �                    �?�㙢�c�?             7@�       �                 �y��?��2(&�?             6@������������������������       �                     &@�       �                 ���?���!pc�?             &@������������������������       �                      @�       �                 p2Ԛ?�����H�?	             "@������������������������       �                     @�       �                 `��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                 �ǋ?П[;U��?             =@�       �                 P�g�?      �?             0@�       �                 ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     �?"pc�
�?             &@�       �                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�θ�?             *@�       �                 @Z�?և���X�?             @������������������������       �                     @�       �                 ���?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                 `.2�?��
ц��?A            @P@�       �                 ����?�g�y��?>             O@�       �                    �?���H.�?2             I@�       �                    �?��S���?-            �F@�       �                     �?�eP*L��?!            �@@�       �                 `dЌ?X�Cc�?             ,@�       �       	             �?�q�q�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 ��f�?      �?              @������������������������       �                     �?������������������������       �                     @�       �                   J�?�����?             3@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?z�G�z�?             .@�       �                 ��3�?؇���X�?             ,@�       �                 �!�?�<ݚ�?	             "@�       �                    �?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?      �?             (@������������������������       �                      @�       �                 ���?ףp=
�?
             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                     �?      �?             (@������������������������       �                     @�       �                 �y�?      �?             @������������������������       �                      @�       �                 @Z�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             8@������������������������       �                      @�       �                    �?"pc�
�?             6@������������������������       �                     @�       �                    �?������?             .@������������������������       �                     �?�       �                 ����?d}h���?             ,@�       �                 pY�?���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	             �?�����H�?	             "@������������������������       �                     @�       �                  ���?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��Q��?             4@�       �                 pg��?      �?              @������������������������       �                     �?�       �                 ����?����X�?             @�       �                    �?r�q��?             @������������������������       �                     @�       �                 `~P�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?r�q��?             (@������������������������       �                     �?�       �                 �:��?�C��2(�?             &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             "@������������������������       �                     @�                       P�c�?&�a2o��?E            @Q@�                       p���?d�;lr�??            �O@�       
      	             �?�d�����?&             C@�       	      
             �?��}*_��?             ;@�       �                 ��8�?�q�q�?             8@�       �                  �Ǩ?�8��8��?             (@������������������������       �        
             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�                          @      �?             (@�       �                 ��a�?����X�?             @������������������������       �                     �?                       �v�?r�q��?             @������������������������       �                     @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?                      �7�?z�G�z�?             @                      ��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@                         @`2U0*��?             9@������������������������       �                     4@                      �-��?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                         �?r�q��?             @������������������������       �                     �?������������������������       �                     @      u                ���?䖏��J�?]           �@                      `p�?ԳC��2�?�             f@������������������������       �                     ?@      J                ��Dz?д>��C�?�             b@      I                   �?�E��ӭ�?6             K@      8                   �?Ȩ�I��?5            �J@      7                   �?���@��?%            �B@      2                P���?4�2%ޑ�?#            �A@                         �?z�G�z�?             >@������������������������       �                     �?      1                p]��?д>��C�?             =@      0                �Єx?�q�q�?             8@       /                   �?�㙢�c�?             7@!      *                ��?z�G�z�?             4@"      )                 DBx?؇���X�?             ,@#      &                @7<x?�<ݚ�?	             "@$      %                �*x?؇���X�?             @������������������������       ��q�q�?             @������������������������       �                     @'      (                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @+      ,                   �?�q�q�?             @������������������������       �                     @-      .                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @3      6                   �?���Q��?             @4      5                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @9      H                P���?      �?             0@:      G                   �?�q�q�?             .@;      F                    �?�eP*L��?             &@<      E                   @���Q��?
             $@=      B                �V�x?�q�q�?	             "@>      A                 ֘�?r�q��?             @?      @                �PHx?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @C      D                p{�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?K      t                   �?L�[2[
�?[            �V@L      k                   �?d1<+�C�?I            @R@M      h                   �?X��Oԣ�?>             O@N      g                �ߵ�?�j��b�?;            �M@O      f                E��?��E�B��?/            �G@P      Y                   �?�q��/��?.             G@Q      T                p��z?`Jj��?             ?@R      S                ��6�?r�q��?             @������������������������       �                     @������������������������       �                     �?U      V                �/��?`2U0*��?             9@������������������������       �                     ,@W      X                 j��?�C��2(�?             &@������������������������       �                     �?������������������������       �        
             $@Z      a                    �?z�G�z�?             .@[      `                   �?����X�?             @\      ]      	             �?r�q��?             @������������������������       �                     @^      _                 ��|?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?b      e                 ""�?      �?              @c      d                `��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     (@i      j                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?l      s                @��?���!pc�?             &@m      n                   �?z�G�z�?
             $@������������������������       �                     �?o      p                   �?�����H�?	             "@������������������������       �                     @q      r                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@v      �                � Q�?"�{	�?�           �z@w      �                   �?X)0���?�            �`@x      y                �?a�?N֩	%��?Y            @V@������������������������       �                     @z      �                P���?X��ʑ��?V            �U@{      �                �x�?h�����?8             L@|      }                �oM�?l��
I��?             ;@������������������������       �                      @~      �                   @�+e�X�?             9@      �                @�X�?�㙢�c�?             7@�      �                   �?����X�?             ,@������������������������       �                     @�      �                s�?      �?              @������������������������       �                      @�      �                ��?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             "@������������������������       �                      @�      �                   �?�f7�z�?             =@�      �                  �?�����H�?	             "@������������������������       �                     �?������������������������       �                      @�      �                  �?�G�z��?             4@�      �                  �?��.k���?             1@������������������������       �                      @�      �                �'t�?��S���?             .@�      �                 �e�?�q�q�?             (@�      �                   �?      �?
             $@������������������������       �                     �?�      �                ��0�?X�<ݚ�?	             "@�      �                ��[�?      �?              @�      �                   �?      �?             @�      �                   @���Q��?             @�      �                �q�?      �?             @������������������������       �                      @�      �                �oM�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                @��?d��0u��?             >@�      �                   �?ףp=
�?
             $@������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?      �?             4@�      �                    �?j���� �?             1@�      �                �q�?�<ݚ�?	             "@�      �      
             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                ��w�?      �?              @�      �                P2`�?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                `o��?�L�lRT�?-            �F@�      �                   �?r٣����?!            �@@������������������������       �                      @�      �                �@�?`�Q��?             9@������������������������       �                      @�      �                 �B�?��+7��?             7@�      �                @y4�?�GN�z�?             6@�      �                �e0�?�t����?             1@�      �                �k�?      �?             0@�      �                 ���?      �?             @������������������������       �                      @������������������������       �                      @�      �                �O��?r�q��?             (@������������������������       �                     @�      �                �ȕ�?�q�q�?             @�      �                P��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                @��?�q�q�?             (@�      �                @x��?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      #                   �?���v{�?'           pr@�      �                 J��?���W�?�            �a@�      �                   @�>����?             ;@�      �                Pn��? �q�q�?             8@�      �                �=��?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     1@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                � W�?�û��|�?s            �\@�      �                p��?"pc�
�?             &@������������������������       �                      @������������������������       �        	             "@�      "                P�s�?$��m��?h             Z@�      �                ���?�q�q�?f            �Y@�      �                ����?���N8�?*             E@�      �                   �?���|���?             6@�      �                 �z�?�z�G��?             4@������������������������       �        	             "@�      �                �q�?�eP*L��?             &@������������������������       �                     @�      �                   �?      �?              @�      �                0���?����X�?             @������������������������       �                      @�      �                    �?���Q��?             @�      �                 x��?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �      
             �?ףp=
�?             4@�      �                ���?�X�<ݺ?             2@�      �                pIz�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@�      �                ����?      �?              @������������������������       �                     �?������������������������       �                     �?�                      �k��?���Q��?<             N@�                      PG��?�����?             3@�                      0�u�?X�<ݚ�?	             "@�                       ��ĩ?և���X�?             @������������������������       �                      @            
             �?���Q��?             @������������������������       �                      @                      �Kŷ?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @            
             �?ףp=
�?
             $@������������������������       �                     @	      
                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                      I9�?���� �?)            �D@������������������������       �                      @      !      	             �?�θ�?'            �C@                         �?��X��?             <@                      2Ѩ?z�G�z�?             4@������������������������       �                     �?                      ���?�S����?             3@                      Х��?$�q-�?             *@                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@                      0��?�q�q�?             @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                       -�?      �?              @                       �2�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@������������������������       �                      @$      %                 ���?��k����?�             c@������������������������       �                     @&      k                �<�?�7�QJW�?�            �b@'      6                ���?�3�o���?�            �b@(      5                �Ѣ?�8��8��?<             N@)      4                 ���?�ݜ�?'            �C@*      3                    �?�KM�]�?&             C@+      ,                ��(�?���y4F�?             3@������������������������       �        
             $@-      .                �\*�?X�<ݚ�?	             "@������������������������       �                      @/      2                ����?����X�?             @0      1                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     3@������������������������       �                     �?������������������������       �                     5@7      f                   �?�����L�?Y            @V@8      O      	             �?�w>�
��?S            �T@9      N                Gm�? �Cc}�?8             L@:      M                ���?"pc�
�?!            �@@;      <                ���?     ��?              @@������������������������       �                     �?=      L                ��Ǹ?��� ��?             ?@>      ?                P�ǲ?ףp=
�?             >@������������������������       �                     ,@@      A                 ��?     ��?             0@������������������������       �                     �?B      K                   �?�r����?             .@C      D                ��4�?�<ݚ�?	             "@������������������������       �                     @E      J                n��?���Q��?             @F      I                   �?�q�q�?             @G      H                ��W�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@P      Q                @Q��?��}*_��?             ;@������������������������       �                      @R      e                   �?`�Q��?             9@S      d                P���?��+7��?             7@T      W                   �?�GN�z�?             6@U      V      
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @X      c                   �?�S����?             3@Y      Z                0��?d}h���?             ,@������������������������       �                     @[      `                ���?�z�G��?
             $@\      _                   �?�q�q�?             @]      ^                `g��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?a      b                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                      @g      h                ��-�?�q�q�?             @������������������������       �                     �?i      j                з~�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?m      �                   �?�Wu�1��?<           �@n      �                   �?Z'8of�?           `q@o      p                p�ҡ?���;�?r            �\@������������������������       �                      @q      z                ��?���X��?p             \@r      y                    �?�����H�?             ;@s      x                ���?�z�G��?
             $@t      w                 �1�?���Q��?             @u      v                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     1@{      �                   �?ҳ�wY;�?U            @U@|      �                   �?և���X�??            �O@}      ~                PUU�?��B����?4             J@������������������������       �                      @      �                   �?      �?2             I@�      �                �l��?p�ݯ��?             3@�      �                �0@�?��
ц��?             *@�      �                �q�?���Q��?
             $@�      �                   @      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                @(��?�P�*�?             ?@�      �                   �?�q�q�?             8@�      �                �tN�?�q�q�?             @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   �?�<ݚ�?             2@�      �                P�c�?$�q-�?             *@������������������������       �                     �?������������������������       �                     (@�      �                p$�?���Q��?             @������������������������       �                      @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                �w�?����X�?             @�      �                   �?r�q��?             @������������������������       �                     @�      �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                �ئ�?"pc�
�?             &@�      �                 	��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                �q�?��2(&�?             6@�      �                   �?      �?             @�      �                 Fж?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�      �                   �?�X�<ݺ?             2@�      �      	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@�      �                 �q�?�p ��?�            �d@�      �                p��?�G�5��?E            @Q@�      �                �'��?4?,R��?$             B@�      �                ����?���Q��?             @������������������������       �                      @�      �                �*�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?`Jj��?             ?@������������������������       �                     2@�      �                �`�?8�Z$���?             *@������������������������       �                     �?�      �                 �q�?�8��8��?             (@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             $@�      �                ���?���|���?!            �@@�      �                �!�?z�G�z�?             .@�      �                ��+�?�z�G��?
             $@�      �                �*��?؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                PUU�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                ��{�?      �?             2@�      �                   �?z�G�z�?
             $@������������������������       �                     �?�      �                @��?�����H�?	             "@�      �                P�%�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   �?      �?              @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                ����?�:nR&y�?_            �W@�      �                   �?      �?@             P@������������������������       �        /            �G@�      �                   �?�t����?             1@������������������������       �        
             $@�      �                    �?����X�?             @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                @���?�חF�P�?             ?@�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @�      �                �RG�?�����H�?             ;@�      �                P_�?     ��?             0@�      �                0���?$�q-�?             *@�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             "@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�      �                   �?�ʱOY��?&           0�@�      k                ����?�2l����?+           �r@�      F      
             �?��#����?�            @l@�      )                �8��?dy�����?�            `c@�                      ��8�?4�M�f��?f            �Y@�                      0��?�q�q�?T             U@�                      �AQ�?�������?D             Q@�      �                `��?b�2�tk�?6             K@�      �                @؀�?�z�G��?
             $@������������������������       �                     @������������������������       �                     @�                      �N�?�X����?,             F@�                      ���?|��?���?             ;@�      �                0���?      �?              @������������������������       �                     @                          �?�q�q�?             @������������������������       �                      @������������������������       �                     �?      
                 �q�?p�ݯ��?             3@                      ����?�q�q�?             (@                         �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @      	                �v!�?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         �?�IєX�?             1@                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@                      ය�?؇���X�?             ,@                         �?$�q-�?             *@                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?            	             �?      �?             0@������������������������       �                     &@                      `�+�?���Q��?             @������������������������       �                     @������������������������       �                      @                          �?�<ݚ�?             2@������������������������       �        	             "@      $                PUU�?X�<ݚ�?	             "@       !                �-I�?z�G�z�?             @������������������������       �                     @"      #                ��!�?      �?              @������������������������       �                     �?������������������������       �                     �?%      (                   �?      �?             @&      '                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @*      ;                   �?�T`�[k�?5            �J@+      4                   �?�S����?&             C@,      3                0?(�?HP�s��?             9@-      2                ���?z�G�z�?
             $@.      1                    �?�����H�?	             "@/      0                ��l�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@5      8                �=��?�	j*D�?             *@6      7                 -��?�����H�?	             "@������������������������       �                     �?������������������������       �                      @9      :                �W��?      �?             @������������������������       �                     @������������������������       �                     �?<      =                �q�?���Q��?             .@������������������������       �                     @>      ?                PUU�?�eP*L��?             &@������������������������       �                      @@      A                   �?X�<ݚ�?	             "@������������������������       �                      @B      C                �uF�?����X�?             @������������������������       �                     @D      E                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?G      j                   �?�ˡ�5��?G            �Q@H      i                0���?V�a�� �?:             M@I      d                 �q�?�*/�8V�?/            �G@J      M                ���?� ��1�?)            �D@K      L                �8��?      �?             0@������������������������       �                     .@������������������������       �                     �?N      O                P���? �o_��?             9@������������������������       �                     �?P      Q                �R�?      �?             8@������������������������       �                     �?R      ]                �;�?��<b���?             7@S      T                   �?�r����?             .@������������������������       �                      @U      \                    �?����X�?             @V      [                   �?      �?             @W      Z      	             �?�q�q�?             @X      Y                `=k�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @^      c                �z��?      �?              @_      `                ����?���Q��?             @������������������������       �                      @a      b                �q�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @e      f                �0%�?�q�q�?             @������������������������       �                     @g      h                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     *@l      y      
             �?��-*��?I            @R@m      r      	             �?�LQ�1	�?             7@n      q                    �?      �?              @o      p                p�R�?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @s      x                   �?z�G�z�?             .@t      u                �8��?      �?              @������������������������       �                     @v      w                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @z      �                ����?���Q��?2             I@{      |                   �?r�q��?             (@������������������������       �                     �?}      ~                Pn��?�C��2(�?             &@������������������������       �        	             "@      �                ���?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                 ��?�\��N��?&             C@������������������������       �                     @�      �                   �?����e��?!            �@@������������������������       �                      @�      �                @q�?f���M�?             ?@�      �                033�?l��
I��?             ;@�      �                 ���?��S���?             .@�      �                �Jk�?���|���?             &@�      �                 ���?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                `(��?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�      �                @8O�?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   �?Hث3���?�           �@�      �                   �?�q�q�?T             U@�      �                p��?���@��?%            �B@�      �      	             �?�	j*D�?             :@�      �                @w\�?��s����?             5@�      �                p̋�?���Q��?             @�      �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                0�b�?      �?             0@������������������������       �                     .@������������������������       �                     �?�      �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�      �                   �?�[�IJ�?/            �G@�      �                   �?�q�q�?             8@�      �                �q�?������?             1@�      �                0���?     ��?             0@�      �                �z��?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �        	             "@������������������������       �                     �?�      �                    �?և���X�?             @������������������������       �                     @�      �                ��8�?      �?             @������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                ��>�?
;&����?             7@������������������������       �                     @�      �                @ �?�G�z��?             4@������������������������       �                     @�      �                Х��?     ��?             0@������������������������       �                      @�      �                ����?      �?             ,@������������������������       �                     @�      �                ����?���|���?             &@������������������������       �                     @�      �                ����?      �?              @�      �                �ǰ�?z�G�z�?             @������������������������       �                     @�      �      
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                PUU�?� ��	��?�           pz@�      �                �ڽ?p�v>��?^            �W@�      �                `K�?�q�q�?             8@������������������������       �                     @�      �                ��t�?�q�q�?             5@�      �                   �?      �?              @������������������������       �                     @�      �                 ��?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                ��I�?��
ц��?             *@�      �                ����?�q�q�?	             "@�      �                @�/�?؇���X�?             @�      �                �f��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�      �                �N.�?z�G�z�?F            �Q@�      �                @q��?(;L]n�?             >@�      �                4��?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@�      �                �^�?�G�z�?(             D@������������������������       �                     @�      �                @�5�?����>�?%            �B@�      �                Ц�?�û��|�?             7@�      �                   @"pc�
�?             &@�      �                 ���?ףp=
�?
             $@�      �                0�G�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                P���?�q�q�?             (@�      �                   �?؇���X�?             @�      �                P�_�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                9��?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                Эm�?@4և���?             ,@������������������������       �                     &@�      �                �E��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                �q�?�^�Q��?I           �t@�      /                   �?�����?+           �r@�                         �?l�;�	�?K            �R@�                      ��8�?��i#[�?*             E@�      �                ��?������?)            �D@������������������������       �                     �?�                       P���?��Q���?(             D@������������������������       �                      @                      ��J�?     ��?              @@                         �?�G�z��?             4@                      �)1�?����X�?             ,@                       �q�?�q�q�?             @������������������������       �                     �?������������������������       �                      @                      ����?"pc�
�?             &@������������������������       �                     @	                      PT�?���Q��?             @
                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                       ��?r�q��?             @                          �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                      �)��?r�q��?             (@                         @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             "@������������������������       �                     �?                      0��?�eP*L��?!            �@@������������������������       �                     @                       ����?l��[B��?             =@                      0��?      �?              @������������������������       �                     @                      ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?!      ,                �@e�?և���X�?             5@"      %      	             �?     ��?             0@#      $                p��?      �?              @������������������������       �                     �?������������������������       �                     @&      +                ����?      �?              @'      (                   @�q�q�?             @������������������������       �                     @)      *                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @-      .                �z�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @0      5                �&��?d}h�m�?�             l@1      2                   �?؇���X�?             @������������������������       �                     @3      4                    �?      �?              @������������������������       �                     �?������������������������       �                     �?6      �                   @�P�*�?�             k@7      8                �q�?o��Ա�?�            `i@������������������������       �                     @9      �                ��?���ׁs�?�             i@:      w                ��?ڇ����?�            @b@;      t                ��_�?�5��?l             [@<      s                `"=�?n�ޢ
�?e            @Y@=      F                �w��?���Q��?_            �W@>      ?                   �?@�0�!��?             1@������������������������       �        	             "@@      E                �|T�?      �?              @A      D                �<�?���Q��?             @B      C                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @G      j                ���?v��:ө�?N            �S@H      c                �^�?     x�?@             P@I      b                `UU�?Tt�ó��?1            �H@J      Y                   �?�lg����?+            �E@K      V                �!��?¦	^_�?             ?@L      U                p�.�?z�G�z�?             9@M      T                {��?�q�q�?             (@N      O                    �?�<ݚ�?	             "@������������������������       �                     �?P      Q                   �?      �?              @������������������������       �                     @R      S                `P��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     *@W      X      	             �?�q�q�?             @������������������������       �                     @������������������������       �                      @Z      a                ��?�q�q�?             (@[      `                 }��?�z�G��?
             $@\      _                ��?      �?             @]      ^                p��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @d      e                p�b�?z�G�z�?             .@������������������������       �                     �?f      g      	             �?؇���X�?             ,@������������������������       �        
             $@h      i                �_��?      �?             @������������������������       �                      @������������������������       �                      @k      n                    �?����X�?             ,@l      m                   �?      �?             @������������������������       �                     @������������������������       �                     �?o      r                �<�?ףp=
�?
             $@p      q                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @u      v                hA=�?؇���X�?             @������������������������       �                     @������������������������       �                     �?x      y                   �?>A�F<�?&             C@������������������������       �                     �?z      {                   �?�MI8d�?%            �B@������������������������       �                     *@|      }                p��?      �?             8@������������������������       �                      @~                      �q�?"pc�
�?             6@������������������������       �                      @�      �                p��?����X�?             ,@������������������������       �                     �?�      �                �G��?�θ�?             *@�      �      	             �?�q�q�?	             "@�      �                ����?      �?              @�      �                    �?؇���X�?             @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                � Q�?      �?6             K@������������������������       �                     @�      �                   �?     ��?0             H@�      �                ��<�?�4�����?             ?@������������������������       �                      @�      �                    �?�c�Α�?             =@�      �                �Ɉ�?X�<ݚ�?	             "@�      �                �8��?z�G�z�?             @������������������������       �                     @�      �                p��?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                05�?      �?             @������������������������       �                     @������������������������       �                     �?�      �                 �q�?R���Q�?             4@�      �                ��[�?�KM�]�?             3@�      �                `�K�?"pc�
�?             &@�      �                `UU�?ףp=
�?
             $@�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                O�?ҳ�wY;�?             1@������������������������       �                     @�      �                ���?d}h���?             ,@�      �                   �?�����H�?	             "@������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                p�g�?���Q��?             @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                ��!�?����X�?             ,@������������������������       �                     @�      �                @&��?X�<ݚ�?	             "@�      �                PAh�?z�G�z�?             @�      �                ��8�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                p���?������?             >@�      �                �q�?d}h���?             <@������������������������       �                     @�      �                `��?����X�?             5@�      �                   �?      �?              @������������������������       �                     @�      �      	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                ���?8�Z$���?             *@������������������������       �                      @�      �                ����?���Q��?             @������������������������       �                      @�      �                   �?�q�q�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      w                �N�?�dG��?�           ؎@�      L                XUU�?������?@            �@�      K                   �?�ՙ/�?�            `b@�      J                �)(y?�%�a�u�?�            �a@�      ?                ��Nc?ꟲ�4��?�            @a@�                      ����?U��K��?y            @^@�      �                   �? �o_��?2             I@������������������������       �                      @�      �                    �?�q�q�?*             E@�      �                @��?���N8�?             5@�      �                 �q?     ��?             0@�      �                �X�?������?             .@�      �                 ��?�q�q�?             (@�      �                   �?�<ݚ�?	             "@�      �                �Z�}?�q�q�?             @������������������������       �                     �?�      �                   @���Q��?             @������������������������       �                     �?�      �                   �?      �?             @������������������������       �                      @�      �                ��`�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                @`ރ?և���X�?             5@�      �                [&�>r�q��?             @������������������������       �                     �?������������������������       �                     @�                         �?��S���?             .@�      �                   @և���X�?             ,@������������������������       �                     �?�      �                ຼ?�n_Y�K�?             *@������������������������       �                     �?�      �                 �q?�q�q�?             (@�      �                ��x�?���Q��?             @�      �                ��d?�q�q�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�                       �!�?����X�?             @������������������������       �                     @                         �?      �?             @                         �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?                      0��%?R_u^|�?G            �Q@                      ��H#?և���X�?             <@	                         �?��
ц��?             *@
                         @�z�G��?
             $@                      P�!?�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �?؇���X�?             @������������������������       �      �?              @������������������������       �                     @������������������������       �                     @                         �?�q�q�?             .@                      �*��?      �?              @                          �?      �?             @������������������������       �                     �?������������������������       �                     @                         �?      �?             @������������������������       �                     �?������������������������       ��q�q�?             @                         �?؇���X�?             @������������������������       �                     @������������������������       �                     �?      <                   �?8�$�>�?+            �E@                         �?V������?%            �B@������������������������       �                     @       ;                   �?�!���?"             A@!      2                @�/?f���M�?             ?@"      1                ��*?���!pc�?             6@#      .                ЉU)?�q�q�?             2@$      -                p�'?d}h���?             ,@%      (                    �?      �?              @&      '                P%O&?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?)      ,                P%O&?z�G�z�?             @*      +                   �?�q�q�?             @������������������������       �      �?              @������������������������       �                     �?������������������������       �                      @������������������������       �                     @/      0                    �?      �?             @������������������������       �      �?              @������������������������       �                      @������������������������       �                     @3      6                P���?X�<ݚ�?	             "@4      5                 wA�?z�G�z�?             @������������������������       ��q�q�?             @������������������������       �                      @7      :                   �?      �?             @8      9                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @=      >                   �?�q�q�?             @������������������������       �                      @������������������������       �                     @@      G                   �?�t����?             1@A      B                   �?@4և���?             ,@������������������������       �        
             $@C      D                    �?      �?             @������������������������       �                      @E      F                ��?      �?              @������������������������       �                     �?������������������������       �                     �?H      I                ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @M      �                0�	�?��]��?�           h�@N      �                   �?�?�P�a�?,           �r@O      �                ����?؍�5���?+           �r@P                       ��?Rԅ5l�?m            @[@Q      j                   �?��|���?X             V@R      ]                   �?ܷ��?��?:             M@S      Z                   �?�}�+r��?&             C@T      Y                   @��?^�k�?#            �A@U      X                ��e�?�8��8��?             (@V      W                ��8�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             $@������������������������       �                     7@[      \                @A �?�q�q�?             @������������������������       �                      @������������������������       �                     �?^      e                   �?z�G�z�?             4@_      d                @�?և���X�?             @`      c                �8��?�q�q�?             @a      b                ��}�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?f      i                ��?$�q-�?             *@g      h                (�q�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@k      z                   �?�������?             >@l      w                0�	�?��2(&�?             6@m      r                ��?ףp=
�?             4@n      o                 �q�?�q�q�?             @������������������������       �                     �?p      q                ���?      �?              @������������������������       �                     �?������������������������       �                     �?s      v                `�2u?�IєX�?             1@t      u                ��Jr?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@x      y                ���?      �?              @������������������������       �                     �?������������������������       �                     �?{      |                    �?      �?              @������������������������       �                     @}      ~                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                �8��?����X�?             5@�      �                ��_r?      �?
             $@������������������������       �                     @�      �                @��?����X�?             @������������������������       �                     @�      �                  �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?�C��2(�?             &@�      �                ��8�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             "@�      �                �q�?�˹�m��?�            �g@�      �                ��[�?̫���/�?�            �a@�      �                   �?��ׄ��?�            `a@�      �                 1��?�E��ӭ�?             2@�      �                �x��?������?             1@�      �                ���?�q�q�?             (@�      �                 �<�?      �?              @������������������������       �                     @������������������������       �                     �?�      �                D)�?      �?             @������������������������       �                      @�      �                `UU�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?0 �����?y            @^@�      �                 ��?�1e�3��?v            �]@�      �                @��? qP��B�?+            �E@������������������������       �        '            �C@�      �                �q=�?      �?             @������������������������       �                     �?������������������������       �                     @�      �                �ئ�?HP�s��?K            �R@�      �                ��R�?     ��?             0@�      �                ��8�?���!pc�?             &@�      �                    �?z�G�z�?
             $@�      �                �@s?      �?             @������������������������       �                     �?�      �                葂�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                �{�p?����˵�?;            �M@�      �                xǡ?      �?             @������������������������       �                     @������������������������       �                     �?�      �                @�?h㱪��?7            �K@������������������������       �                      @@�      �                `�ک?���}<S�?             7@�      �                   @����X�?             @�      �                   �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@�      �                P(��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                 �	�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        0             H@������������������������       �                     �?�      �                �66�?4�2%ޑ�?�           x@�      �                   �?|��?���?             ;@�      �                ����?r�q��?             8@�      �                @�h�?�ՙ/�?             5@�      �                �{B�?      �?             ,@�      �      	             �?���|���?             &@�      �                ���?؇���X�?             @������������������������       �                     �?������������������������       �                     @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?؇���X�?             @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      v                PUU�?,m�)6��?f           `v@�      ;                   �?4��s?D�?J           �t@�      ,                ���?t�R2��?�            �k@�      	                   �?fv�S��?�            �d@�      �                ��'�?R�(CW�?R            �T@�      �                   �?�q�q�?             (@������������������������       �                     @�      �                Po�?�<ݚ�?	             "@�      �                   �?      �?              @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�                      p��?(N:!���?F            �Q@�      �      	             �?�θV�?E            @Q@�      �                   �?���N8�?*             E@������������������������       �                     7@�      �                @���?�KM�]�?             3@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   @�IєX�?             1@������������������������       �                     *@�      �                ����?      �?             @������������������������       �                      @�      �                �a��?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   @�+$�jP�?             ;@�      �                   �?�����H�?             2@�      �                �q�?      �?             0@�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@�      �                 =�?      �?              @������������������������       �                     �?������������������������       �                     �?                       �w�?�q�q�?	             "@������������������������       �                     �?                      P�E�?      �?              @                      �$A�?؇���X�?             @������������������������       �                     @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?
      %                ��8�?��p �?R            �T@                      ��8�?     x�?@             P@                         �?4�2%ޑ�?#            �A@                      �:B�?�8��8��?             8@������������������������       �                     5@                      ��?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �?�eP*L��?             &@������������������������       �                     @                      ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @      "                �V��?l��[B��?             =@                         @�z�G��?             4@                      ����?     ��?             0@������������������������       �                     @                         �?�q�q�?	             "@������������������������       �                     @                         �?���Q��?             @������������������������       �                     @������������������������       �                      @       !                   �?      �?             @������������������������       �                     @������������������������       �                     �?#      $                P�&�?�����H�?	             "@������������������������       �                      @������������������������       �                     �?&      +                 Y��?�����H�?             2@'      (      
             �?�IєX�?             1@������������������������       �                     .@)      *                ��\�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?-      :                    �? ,��-�?;            �M@.      /                   �?      �?              @@������������������������       �                     *@0      1                �^4�?���y4F�?             3@������������������������       �                     �?2      9                �S��?r�q��?             2@3      8                   �?�t����?             1@4      5      	             �?�q�q�?             @������������������������       �                     @6      7                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                     ;@<      =                ����?xZ�l ��?k            �Z@������������������������       �                      @>      m                   �?����X�?i            @Z@?      R                   �?>���Rp�?W            �U@@      K                �<t�?ZՏ�m|�?1            �H@A      H                   �?��(\���?(             D@B      C                   �?��?^�k�?#            �A@������������������������       �                     8@D      E                   �?�C��2(�?             &@������������������������       �                     @F      G                p��?      �?             @������������������������       �                     �?������������������������       �                     @I      J                @_r�?���Q��?             @������������������������       �                      @������������������������       �                     @L      Q                   �?X�<ݚ�?	             "@M      P                �X��?r�q��?             @N      O                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @S      V                 ���?P����?&             C@T      U                �� �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @W      X                p	��?���!pc�?!            �@@������������������������       �                     �?Y      `                   �?      �?              @@Z      _                ���?�t����?             1@[      \                �8��?���Q��?             @������������������������       �                      @]      ^                0�	�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@a      f                �2�?���Q��?             .@b      e                   �?�q�q�?             @c      d                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?g      h                   �?�<ݚ�?	             "@������������������������       �                     �?i      j                �#��?      �?              @������������������������       �                     @k      l                    �?      �?              @������������������������       �                     �?������������������������       �                     �?n      o                0���?      �?             2@������������������������       �                     @p      q                   �?X�Cc�?             ,@������������������������       �                     @r      u                �k��?X�<ݚ�?	             "@s      t                 �յ?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     <@x      �                ��J�?b�MKm�?�            `c@y      �                �rv�?����5�?=            �N@z      �                   �?�E��ӭ�?6             K@{      �                �~��?��S���?             .@|                      ����?      �?              @}      ~                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   @؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                ���?:�&���?'            �C@�      �                ��?ҳ�wY;�?             1@�      �                ����?������?             .@������������������������       �                     @�      �                ��8�?      �?              @������������������������       �                      @�      �                   �?�q�q�?             @�      �                p��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�      �                    �?���7�?             6@������������������������       �                     .@�      �                @A*�?؇���X�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                �8��?����X�?             @������������������������       �                      @������������������������       �                     @�      �                 R��?@�҇��?^            �W@�      �                �ۋ�?���*~�?Y            @V@�      �                �q�?����X�?8             L@�      �                0=P�?�q�q��?0             H@�      �                   �?��S�ۿ?             .@������������������������       �                     &@�      �                0)��?      �?             @������������������������       �                     �?������������������������       �                     @�      �                ���?:ɨ��?!            �@@�      �                �q�?և���X�?             5@�      �                   @�t����?             1@�      �      
             �?      �?             0@�      �                   �?���Q��?
             $@������������������������       �                     @�      �                p��?և���X�?             @������������������������       �                      @�      �                   �?���Q��?             @������������������������       �                      @�      �                 ~��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?�8��8��?             (@������������������������       �        	             "@�      �      	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                P��?      �?              @������������������������       �                     @�      �                O\�?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   �?�C��2(�?!            �@@�      �                ���?      �?              @������������������������       �                     @�      �                ��X�?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?`2U0*��?             9@�      �      	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�      �                 q��?z�G�z�?             @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                P�?�M���?�	           �@�      �                   �?،(��?�           �@�      @                   �?x��ėb�?w           ��@�                      �ae�?P;ߣ	H�?|           ��@�      �                 �Fa? �t��̮?�           0|@�      �                �J_?z�G�z�?
             $@�      �                   �?�����H�?	             "@�      �                XUU�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?P����?�           �{@�      �                ����?�U�=���?B            �P@������������������������       �                     �?�      �                `�ת?����?A            @P@�      �                �iF�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?P���Q�?<             N@������������������������       �                     ;@�      �                �A�?�C��2(�?!            �@@�      �                ��N�?��2(&�?             6@�      �                   �?�����?             5@�      �                p��?�}�+r��?             3@������������������������       �                     0@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�                         @�v¢?w           pw@�      �                   �? f^8���?�            �i@�      �                   �?PA��ڡ?�             e@�      �                 ��?XB���?W            �U@������������������������       �        !            �@@�      �                �*��?�X�<ݺ?6             K@������������������������       �                     �?�      �                ���?�&=�w��?5            �J@�      �                �|��?@4և���?             <@�      �                �q�? 7���B�?             ;@������������������������       �                     5@�      �                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     9@������������������������       �        R            �T@                           �?�L���?%            �B@������������������������       �                     1@                         �?R���Q�?             4@                         �?���!pc�?             &@������������������������       �                     �?                      PUU�?z�G�z�?
             $@������������������������       �                     @      
                   �?���Q��?             @      	                �1��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        	             "@                      �Fj�?@�����?�             e@                      ����?�IєX�?             1@������������������������       �                     0@������������������������       �                     �?������������������������       �        �             c@                      ���?�L���?�             g@                      ���?�	j*D�?             *@                      p�Ǽ?"pc�
�?             &@������������������������       �                     �?                         �?ףp=
�?
             $@������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @      5                �8��?�Ts�k��?�            �e@      4                Ё��?t�U����?C            �P@      1                ����?��IF�E�?B            �P@      (                   @�8��8��?<             N@       %                �[�?`�q�0ܴ?/            �G@!      $                P���?��Y��]�?)            �D@"      #                `���?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     =@&      '                0j��?r�q��?             @������������������������       �                     �?������������������������       �                     @)      ,                   �?�θ�?             *@*      +                @�2�?�q�q�?             @������������������������       �                      @������������������������       �                     �?-      .                ��?ףp=
�?
             $@������������������������       �                     @/      0                �p�?�q�q�?             @������������������������       �                     �?������������������������       �                      @2      3                0t�?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?6      7                �$��?��?^�k�?i            @Z@������������������������       �        V            �U@8      9                   �?�S����?             3@������������������������       �                     (@:      ;                ��E�?և���X�?             @������������������������       �                      @<      ?                �q�?z�G�z�?             @=      >                ��5�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @A      P                �	��?�vps�?�            `o@B      C                @kg�?�q�q�?             5@������������������������       �                      @D      M                @#�?�d�����?             3@E      J                ;x�?     ��?             0@F      I                �RG�?ףp=
�?
             $@G      H                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @K      L                �n��?�q�q�?             @������������������������       �                      @������������������������       �                     @N      O                �q�?�q�q�?             @������������������������       �                      @������������������������       �                     �?Q      Z                �t:�?���AY5�?�            �l@R      S                �0@�?�g�y��?>             O@������������������������       �        6             K@T      U                �o�?      �?              @������������������������       �                     �?V      W                   �?؇���X�?             @������������������������       �                     @X      Y                   �?      �?              @������������������������       �                     �?������������������������       �                     �?[      ^                �̱�?�X�C�?�             e@\      ]                0��?      �?             @������������������������       �                     �?������������������������       �                     @_      ~                `�b�?�p ��?�            �d@`      o      	             �?d��0u��?<             N@a      n                �U�?�t����?"             A@b      e                `UU�?�C��2(�?!            �@@c      d                   �?      �?              @������������������������       �                     �?������������������������       �                     �?f      g                �ri�?`Jj��?             ?@������������������������       �                     4@h      m                   �?"pc�
�?             &@i      j                `�A�?ףp=
�?
             $@������������������������       �                     @k      l                `�t�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?p      u                ��#�?$��m��?             :@q      t                 �z�?և���X�?             @r      s      
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @v      w                ����?�d�����?             3@������������������������       �                     @x      y                P��?�q�q�?             (@������������������������       �                     @z      }                   �?����X�?             @{      |                   @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?      �                �q
�?,�T�6�?h             Z@������������������������       �                     �?�      �                `kB�?p���p�?g            �Y@������������������������       �                     <@�      �                Ж��?�r����?K            �R@������������������������       �                     �?�      �                   @��(�2Y�?J            �R@�      �                �ئ�?�θV�?E            @Q@�      �                P8O�?���c���?4             J@�      �                ��]�?�t����?3            �I@�      �                �MF�?�:�^���?-            �F@�      �                �PT�?�7��?'            �C@�      �                 �=�?�r����?             .@�      �                p��?@4և���?             ,@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     �?������������������������       �                     8@�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     @�      �                �q��?�q�q�?             @������������������������       �                     �?�      �                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     1@�      �                   �?���Q��?             @������������������������       �                     @������������������������       �                      @�      �                0���? @ެ[�?           @�@�      �                ���? D�R��?3           ��@�      �                PHy�?����3�?1           ��@�      �                �q�?�����?�            �@�      �                PUU�?��Vl��?�           `{@�      �                ����?�:!�g��?X           �u@������������������������       �        �             g@�      �                P���?Уp=
ע?�             d@�      �                ����?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                �?�Fǌ��?�            �c@�      �                0X~�?r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   �? i�*$Ŋ?�             c@�      �                ����?г�wY;�?"             A@�      �                `��?$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     5@������������������������       �        v            �]@�      �                    �?`�q�0ܴ?^            �W@������������������������       �        .             G@�      �                �B#�?�8��8��?0             H@�      �                �&��?���Q��?             @������������������������       �                      @�      �                �S��?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                �q�? �#�Ѵ�?+            �E@�      �                ��8�?�C��2(�?             6@������������������������       �                     &@�      �      
             �?"pc�
�?             &@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                �"��?�����H�?	             "@�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     5@�      �                   �? ��e{?*           �r@�      �                p��?XB���?             =@������������������������       �                     ;@�      �      
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                   �p@�      �                 ��? 7���B�?Q            @T@������������������������       �                     �?�      �      	             �?�(\����?P             T@�      �                �"X�?�t����?             1@������������������������       �                     �?�      �      
             �?      �?             0@�      �                ��?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �        ?            �O@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        �            �k@�      z                   �?r�q��?p           ��@�      u                �N�?�+e�X�?E           Pt@�      t                PUU�?�t����??           �s@�                      ���?Z�/�j��?*           �r@�      �                `��?������?[            �V@�      �                ���?�t����?             1@�      �                   �?z�G�z�?             .@������������������������       �        	             "@�      �                   �?      �?             @������������������������       �                      @�      �                `�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�                      �8��?$G$n��?J            �R@�                         �? ���g=�?E            @Q@�                      `���?ZՏ�m|�?1            �H@�                         �?8��8���?0             H@�      �                   �?tk~X��?$             B@�      �                P��?�q�q�?             (@�      �      	             �?և���X�?             @�      �                ��_�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   �?      �?             8@������������������������       �        	             "@�      �                �q�?z�G�z�?             .@������������������������       �                     @�                          �?�q�q�?	             "@������������������������       �                     @                      �B��?      �?             @                      ��8�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                     �?������������������������       �                     4@	      
      
             �?���Q��?             @������������������������       �                      @������������������������       �                     @      U                `q'�?�m淣�?�            �i@      8                p��?�X���?�            �`@      !      
             �?���mC�?U            @U@                          �?r�q��?             8@                      mQ�?�G�z��?             4@                       ��?�n_Y�K�?             *@������������������������       �                      @                      �8��?���!pc�?             &@                       �G�?      �?             @                      �{�?      �?             @            	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                          �?؇���X�?             @������������������������       �                     @                      `��?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @"      #                p��?`��:�?=            �N@������������������������       �                     ,@$      %                p���?�*/�8V�?/            �G@������������������������       �                      @&      -      	             �?�<ݚ�?-            �F@'      (                ph��?ҳ�wY;�?             1@������������������������       �                     @)      *                �e�?d}h���?             ,@������������������������       �                      @+      ,                    �?      �?             @������������������������       �                     @������������������������       �                     @.      1                   �?؇���X�?             <@/      0                   �?��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@2      7                @?��?�θ�?             *@3      6                ����?      �?             @4      5                �M�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @9      H                   �?JJ����?/            �G@:      ?                   �?�û��|�?             7@;      <                ����?�����H�?	             "@������������������������       �                     @=      >                 ���?      �?              @������������������������       �                     �?������������������������       �                     �?@      A                   �?և���X�?             ,@������������������������       �                     @B      C                ����?���Q��?
             $@������������������������       �                     @D      G                ��k�?և���X�?             @E      F                ���?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @I      T                ����?�q�q�?             8@J      K                 ���?���!pc�?             6@������������������������       �                     @L      M                Pc�?      �?             0@������������������������       �                     @N      O                `UU�?�θ�?             *@������������������������       �                     @P      S                 �1�?և���X�?             @Q      R                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @V      m                `4O�?��n�?K            �R@W      l                   �?؇���X�??            �O@X      Y                `�m�?�θ�?'            �C@������������������������       �                     �?Z      k                   �?���y4F�?&             C@[      \                ��I�?`�Q��?             9@������������������������       �                     @]      h                   �?X�<ݚ�?             2@^      _                   �?      �?             (@������������������������       �                     �?`      g                �%�?"pc�
�?             &@a      f                �V��?�q�q�?             @b      c                �Ջ�?z�G�z�?             @������������������������       �                     @d      e                 ���?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @i      j                @Ӭ�?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     8@n      o                Pq��?�q�q�?             (@������������������������       �                     @p      s                ����?      �?              @q      r      	             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     5@v      y                   �?�q�q�?             @w      x                �mu�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @{      �                ��,�?���}<S�?+           �r@|                      p۶�?���Q��?             @}      ~                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                p��?��v�u�?&           `r@�      �                `���?pb����?�             g@�      �                 �J�?p�qG�?`             X@�      �                ���?r�q��?             8@�      �                �rv�?�LQ�1	�?             7@�      �                p2��?�C��2(�?             6@�      �                ��?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     0@������������������������       �                     �?������������������������       �                     �?�      �                �_��?�k~X��?H             R@�      �                 �p�?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �        9            �L@�      �                p�#�?NKF����?Y            @V@�      �                �8��?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                ��8�?0,Tg��?T             U@�      �                0��?����X�?             <@�      �                   �?"pc�
�?             6@������������������������       �        	             "@�      �                0���?�	j*D�?             *@�      �                   �?      �?              @������������������������       �                      @�      �                 ��?�q�q�?             @������������������������       �                     @�      �                �v4�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                 S�?�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                   �?4և����?8             L@�      �                 .�?     ��?             0@�      �                p��?�r����?             .@�      �                ��8�?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             $@������������������������       �                     �?�      �                0Io�?P���Q�?(             D@������������������������       �                     6@�      �                ����?�����H�?             2@������������������������       �                     �?�      �                �q�?�IєX�?             1@�      �                гv�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@�      �                 �>�?��wڝ�?m            @[@�      �                P�?�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?������������������������       �        Z            �V@��      �t�b�values�hhK ��h��R�(KM�KK��hx�B��       *�@     `�@     ��@     ��@      �@     ��@      w@     �@     �i@      i@      c@      g@     �O@     �Z@     �H@     �P@     �H@      M@     �G@     �G@      D@      G@     �A@     �F@      9@      7@      8@      0@      .@      @      &@      @      &@      @      @       @               @      @               @      �?      @              �?      �?              �?      �?                       @      @              "@      &@      @      @      @      @       @      @              �?       @      @      �?              �?      @      �?      �?              �?      �?                       @      �?                      @      @      @      �?      @      �?                      @      @      �?       @      �?       @                      �?      @              �?      @              @      �?              $@      6@      @      5@      @      3@              &@      @       @      @      @       @      @       @      �?              �?       @                      @      �?                      @      @       @      �?       @              �?      �?      �?      �?                      �?       @              @      �?              �?      @              @      �?              �?      @              @      �?      @              �?      �?      �?                      �?       @      &@       @      @      �?      @              @      �?       @      �?                       @      �?                      @               @      ,@      D@      @      A@      �?      .@              *@      �?       @               @      �?              @      3@      @      2@      �?      &@      �?       @               @      �?                      "@      @      @       @              �?      @      �?      �?      �?                      �?              @       @      �?              �?       @              @      @      @              @      @      �?      @              @      �?      �?              �?      �?               @             �V@     �S@     �V@      R@     �T@     �M@     @P@     �J@     �A@      2@      3@      @      3@      @      3@      @      &@               @      @               @       @      �?      @               @      �?       @                      �?              �?              �?      0@      *@      @      $@      @      �?              �?      @               @      "@       @       @       @                       @              @      $@      @      @      @      @              �?      @              @      �?              @              >@     �A@      >@      @@      5@      =@      5@      8@      2@      .@      @      "@      @       @      @              �?       @      �?                       @      �?      @      �?                      @      *@      @      �?      @              @      �?              (@      @      (@       @      @       @      @      �?      @               @      �?       @                      �?              �?      @                      �?      @      "@       @              �?      "@              @      �?       @      �?                       @              @      "@      @      @              @      @               @      @      �?      @                      �?              @      2@      @               @      2@      @      @              &@      @              �?      &@      @      @       @       @              �?       @      �?                       @       @      �?      @              �?      �?              �?      �?              @      *@      @      @              �?      @       @      @      �?      @               @      �?       @                      �?              �?       @      $@      �?              �?      $@      �?      �?              �?      �?                      "@              @     �J@      0@      J@      &@      <@      $@      1@      $@      1@      @      &@      �?      $@              �?      �?              �?      �?              @      @       @      @      �?              �?      @              @      �?      �?      �?                      �?      @      �?      �?      �?      �?                      �?      @                      @      &@              8@      �?      4@              @      �?      @                      �?      �?      @      �?                      @     �d@     �{@      9@     �b@              ?@      9@      ^@      .@     �C@      ,@     �C@       @      =@       @      ;@      @      8@      �?              @      8@      @      3@      @      3@      @      0@       @      (@       @      @      �?      @      �?       @              @      �?      �?      �?                      �?              @       @      @              @       @      �?              �?       @                      @      �?                      @       @      @       @      �?              �?       @                       @               @      @      $@      @      $@      @      @      @      @      @      @      �?      @      �?       @               @      �?                      @       @      �?       @                      �?      �?              �?                      @      �?              �?              $@     @T@      $@     �O@      @     �K@      @     �J@      @     �D@      @     �D@       @      =@      �?      @              @      �?              �?      8@              ,@      �?      $@      �?                      $@      @      (@       @      @      �?      @              @      �?      �?      �?                      �?      �?              �?      @      �?       @               @      �?                      @      �?                      (@      �?       @               @      �?              @       @       @       @      �?              �?       @              @      �?       @               @      �?              �?                      2@     `a@      r@     �O@     �Q@     �G@      E@      @              F@      E@      9@      ?@       @      3@       @              @      3@      @      3@      @      $@              @      @      @               @      @       @      @                       @              "@       @              1@      (@       @      �?              �?       @              "@      &@      "@       @       @              @       @      @      @      @      @      �?              @      @      @      @      @      @      @       @      @      �?       @              �?      �?              �?      �?                      �?              �?               @      �?               @                      @              @      3@      &@      "@      �?       @              �?      �?              �?      �?              $@      $@      $@      @      @       @       @       @       @                       @      @              @      @      @       @               @      @                      @              @      0@      =@       @      9@               @       @      1@       @              @      1@      @      1@      @      (@      @      (@       @       @               @       @               @      $@              @       @      @       @      �?       @                      �?              @      �?                      @      �?               @      @       @      @       @                      @      @              S@     `k@     �G@     �W@       @      9@      �?      7@      �?      @              @      �?                      1@      �?       @      �?                       @     �F@     �Q@      "@       @               @      "@              B@      Q@      A@      Q@      $@      @@       @      ,@      @      ,@              "@      @      @      @              @      @       @      @               @       @      @       @      �?       @                      �?               @      �?               @               @      2@      �?      1@      �?      @              @      �?                      *@      �?      �?              �?      �?              8@      B@      *@      @      @      @      @      @       @               @      @               @       @      �?       @                      �?               @      "@      �?      @               @      �?       @                      �?      &@      >@       @              "@      >@      "@      3@      @      0@      �?              @      0@      �?      (@      �?      �?              �?      �?                      &@       @      @       @      �?              �?       @                      @      @      @      �?      @      �?                      @      @                      &@       @              =@      _@      @              :@      _@      9@      _@      @     �K@      @      A@      @      A@      @      .@              $@      @      @       @               @      @       @      �?              �?       @                      @              3@      �?                      5@      4@     @Q@      0@     �P@      @      I@      @      ;@      @      ;@      �?              @      ;@      @      ;@              ,@      @      *@      �?               @      *@       @      @              @       @      @       @      �?      �?      �?              �?      �?              �?                       @              @      �?              �?                      7@      $@      1@       @               @      1@      @      1@      @      1@       @      �?              �?       @              @      0@      @      &@              @      @      @       @      �?      �?      �?      �?                      �?      �?              �?      @      �?                      @              @      �?               @              @       @              �?      @      �?      @                      �?      �?             p�@     �z@     `k@     �M@     �S@     �A@               @     �S@     �@@      8@      @      @      @       @      @       @      �?       @                      �?               @      @              1@             �K@      >@      B@      ;@      ;@      9@       @              9@      9@      @      (@      @      @      @      @       @      @              @       @               @              @                      @      2@      *@      0@       @       @      @       @      �?              �?       @                      @      ,@      @      (@      �?              �?      (@               @      @               @       @      �?              �?       @               @      @      �?      @              @      �?      �?              �?      �?              �?              "@       @      �?       @      �?                       @       @              3@      @       @       @       @      �?       @                      �?              �?      1@      �?       @      �?              �?       @              .@             �a@      8@      J@      1@      ?@      @       @      @               @       @      �?       @                      �?      =@       @      2@              &@       @              �?      &@      �?      �?      �?      �?                      �?      $@              5@      (@      (@      @      @      @      @      �?      @                      �?      �?       @      �?                       @      @              "@      "@       @       @      �?              �?       @      �?       @               @      �?                      @      @      �?       @      �?       @                      �?      @              V@      @      O@       @     �G@              .@       @      $@              @       @      �?       @      �?                       @      @              :@      @       @       @       @                       @      8@      @      *@      @      (@      �?      @      �?      @                      �?      "@              �?       @      �?                       @      &@             0{@     0w@     �g@     �[@      c@     @R@     �W@     �N@     �J@     �H@     �H@     �A@     �A@     �@@     �@@      5@      @      @      @                      @      >@      ,@      ,@      *@      @      �?      @               @      �?       @                      �?      @      (@      @      @      �?      @      �?                      @      @      �?              �?      @                      @      0@      �?       @      �?       @                      �?      ,@               @      (@      �?      (@      �?      �?      �?                      �?              &@      �?              ,@       @      &@              @       @      @                       @      @      ,@              "@      @      @      �?      @              @      �?      �?      �?                      �?      @      �?      �?      �?              �?      �?               @             �D@      (@      @@      @      7@       @       @       @       @      �?       @      �?              �?       @              @                      �?      .@              "@      @       @      �?              �?       @              �?      @              @      �?              "@      @      @              @      @               @      @      @               @      @       @      @              �?       @               @      �?             �M@      (@      G@      (@     �A@      (@     �@@       @      .@      �?      .@                      �?      2@      @              �?      2@      @              �?      2@      @      *@       @       @              @       @       @       @       @      �?      �?      �?              �?      �?              �?                      �?      @              @      @       @      @               @       @      �?       @                      �?      @               @      @              @       @      �?              �?       @              &@              *@             �A@      C@      .@       @      @      @      @       @               @      @                      @      (@      @      @      @      @              �?      @              @      �?              @              4@      >@       @      $@      �?              �?      $@              "@      �?      �?      �?                      �?      2@      4@      @              *@      4@       @              &@      4@       @      3@      @       @      @      @      �?      @              @      �?              @                      @      �?      &@      �?                      &@      @      �?      @                      �?     �n@     @p@      L@      <@      =@       @      2@       @      1@      @       @      @       @      �?              �?       @                       @      .@      �?      .@                      �?      �?      @              @      �?              &@              ;@      4@      0@       @      *@      @      *@      @      @      @      @                      @      "@                      �?      @      @              @      @      �?       @              �?      �?              �?      �?              &@      (@              @      &@      "@      @              @      "@               @      @      @      @              @      @              @      @      @      @      �?      @              �?      �?      �?                      �?              @     �g@      m@      <@     �P@      ,@      $@              @      ,@      @      @      �?      @              �?      �?              �?      �?              @      @      @      @      �?      @      �?      �?              �?      �?                      @       @              @              ,@      L@      �?      =@      �?      @              @      �?                      9@      *@      ;@      @              $@      ;@      "@      ,@       @      "@      �?      "@      �?      �?      �?                      �?               @      �?              @      @      @      �?      �?      �?      �?                      �?      @              �?      @      �?                      @      �?      *@              &@      �?       @               @      �?             `d@     �d@     �a@     �c@      F@      ?@      =@      *@      =@      (@              �?      =@      &@       @              5@      &@      &@      "@      $@      @      �?       @      �?                       @      "@       @      @              @       @      �?       @      �?                       @       @              �?      @      �?      �?              �?      �?                      @      $@       @      �?       @               @      �?              "@                      �?      .@      2@              @      .@      ,@      @       @      @              �?       @               @      �?              "@      (@      @      &@      �?      @      �?                      @      @      @      @       @      @              �?       @               @      �?                       @      @      �?              �?      @             @X@     �_@      @      �?      @              �?      �?              �?      �?             �V@     �_@     @T@     �^@      @             �S@     �^@     �I@     �W@      F@      P@      C@     �O@      C@     �L@      @      ,@              "@      @      @      @       @      �?       @      �?                       @       @                      @     �A@     �E@      9@     �C@      6@      ;@      0@      ;@      "@      6@      @      4@      @      @       @      @      �?              �?      @              @      �?      �?      �?                      �?      @                      *@      @       @      @                       @      @      @      @      @      �?      @      �?      �?      �?                      �?               @      @                       @      @              @      (@      �?               @      (@              $@       @       @       @                       @      $@      @      �?      @              @      �?              "@      �?      �?      �?      �?                      �?       @                      @      @      �?      @                      �?      @      ?@      �?              @      ?@              *@      @      2@       @              @      2@               @      @      $@      �?              @      $@      @      @       @      @      �?      @      �?       @               @      �?                      @      �?              �?                      @      ;@      ;@      @              5@      ;@      $@      5@       @               @      5@      @      @      @      �?      @              �?      �?              �?      �?              �?      @              @      �?              @      1@       @      1@       @      "@      �?      "@      �?       @               @      �?                      @      �?                       @      �?              &@      @              @      &@      @       @      �?      @               @      �?              �?       @              @       @      �?       @               @      �?               @              $@      @      @              @      @      �?      @      �?      �?              �?      �?                      @      @              6@       @      6@      @      @              .@      @      @      @      @              �?      @      �?                      @      &@       @       @              @       @       @              �?       @      �?      �?      �?                      �?              �?               @     @�@     `n@     h�@     `f@     �V@      L@     �V@     �I@     �V@     �G@      S@     �F@      B@      ,@       @              <@      ,@      0@      @      &@      @      &@      @       @      @      @       @      @       @      �?              @       @              �?      @      �?       @              �?      �?              �?      �?              @              �?       @               @      �?              @                      �?      @              (@      "@      @      �?              �?      @              @       @      @       @      �?              @       @              �?      @      @      @       @      �?       @      �?      �?              �?      �?                      �?       @               @      @              @       @       @       @      �?      �?      �?      �?                      �?      �?              D@      ?@      (@      0@      @      @      @      @      �?       @      �?                       @      @      �?      �?      �?      @                      @      @      $@      @      @      �?      @      �?                      @      @      �?      �?               @      �?      �?      @              @      �?              <@      .@      :@      &@      @              7@      &@      4@      &@      0@      @      (@      @      &@      @      @      @      �?       @      �?      �?              �?      @      �?       @      �?      �?      �?      �?               @              @              �?      @      �?      �?               @      @              @      @      �?      @      �?       @               @      @      �?      �?      �?      �?                      �?       @              @               @      @       @                      @      .@       @      *@      �?      $@              @      �?       @              �?      �?      �?                      �?       @      �?              �?       @                      @              @     ��@     �^@     �p@     �A@     �p@      A@     �V@      3@     �R@      *@      J@      @      B@       @      A@      �?      &@      �?      �?      �?              �?      �?              $@              7@               @      �?       @                      �?      0@      @      @      @      @       @      �?       @               @      �?              @                      �?      (@      �?      �?      �?      �?                      �?      &@              7@      @      3@      @      2@       @       @      �?      �?              �?      �?              �?      �?              0@      �?      @      �?      @                      �?      (@              �?      �?      �?                      �?      @      @              @      @      �?              �?      @              .@      @      @      @      @               @      @              @       @      �?       @                      �?      $@      �?      �?      �?      �?                      �?      "@             �e@      .@     �_@      .@     �_@      *@      *@      @      *@      @       @      @      @      �?      @                      �?      �?      @               @      �?      �?              �?      �?              @                      �?     @\@       @     �[@      @      E@      �?     �C@              @      �?              �?      @             @Q@      @      *@      @       @      @       @       @       @       @      �?              �?       @               @      �?              @                      �?      @              L@      @      @      �?      @                      �?     �J@       @      @@              5@       @      @       @      @      �?      @                      �?              �?      0@               @      �?       @                      �?      �?       @               @      �?              H@                      �?     �r@      V@      *@      ,@      *@      &@      *@       @      @      @      @      @      @      �?              �?      @              �?      @              @      �?                      @      @      �?      @              �?      �?      �?                      �?              @              @     �q@     �R@      p@     �R@     �f@      E@     �_@      C@     @Q@      *@      @      @              @      @       @      @      �?      �?      �?      �?                      �?      @                      �?      O@       @      O@      @      D@       @      7@              1@       @      �?      �?      �?                      �?      0@      �?      *@              @      �?       @              �?      �?              �?      �?              6@      @      0@       @      .@      �?       @      �?       @                      �?      *@              �?      �?      �?                      �?      @      @              �?      @       @      @      �?      @              �?      �?              �?      �?                      �?              �?     �L@      9@     �D@      7@      ;@       @      6@       @      5@              �?       @      �?                       @      @      @      @              �?      @      �?                      @      ,@      .@      @      ,@      @      *@              @      @      @              @      @       @      @                       @      @      �?      @                      �?       @      �?       @                      �?      0@       @      0@      �?      .@              �?      �?      �?                      �?              �?     �K@      @      <@      @      *@              .@      @              �?      .@      @      .@       @      @       @      @              �?       @               @      �?              &@                      �?      ;@             �R@      @@               @     �R@      >@     �P@      5@     �D@       @     �B@      @      A@      �?      8@              $@      �?      @              @      �?              �?      @              @       @               @      @              @      @      �?      @      �?      �?      �?                      �?              @      @              9@      *@      �?      @      �?                      @      8@      "@              �?      8@       @      .@       @      @       @       @              �?       @               @      �?              (@              "@      @       @      @      �?      @      �?                      @      �?              @       @              �?      @      �?      @              �?      �?      �?                      �?      "@      "@              @      "@      @      @              @      @      @      �?              �?      @                      @      <@             �V@      P@      4@     �D@      .@     �C@       @      @       @      @       @      �?              �?       @                      @      @      �?      @                      �?      @      @@      @      &@      @      &@              @      @      @       @               @      @       @      �?              �?       @                      @       @              �?      5@              .@      �?      @      �?      �?              �?      �?                      @      @       @               @      @             �Q@      7@     �Q@      3@      D@      0@     �B@      &@      ,@      �?      &@              @      �?              �?      @              7@      $@      (@      "@      (@      @      (@      @      @      @      @              @      @               @      @       @       @              �?       @      �?                       @      @                      �?              @      &@      �?      "@               @      �?              �?       @              @      @              @      @      �?      @                      �?      >@      @      @       @      @              �?       @      �?                       @      8@      �?      @      �?              �?      @              4@              �?      @              @      �?      �?              �?      �?             ��@     �f@     �@     @S@     ��@     @P@     ��@      =@     P{@      ,@       @       @       @      �?      �?      �?      �?                      �?      @                      �?     �z@      (@     �N@      @              �?     �N@      @      @      �?      @                      �?     �L@      @      ;@              >@      @      3@      @      3@       @      2@      �?      0@               @      �?              �?       @              �?      �?              �?      �?                      �?      &@              w@      @      i@      @     �d@      @      U@      @     �@@             �I@      @              �?     �I@       @      :@       @      :@      �?      5@              @      �?              �?      @                      �?      9@             �T@              A@      @      1@              1@      @       @      @              �?       @       @      @              @       @      �?       @      �?                       @       @              "@              e@      �?      0@      �?      0@                      �?      c@             @e@      .@      "@      @      "@       @              �?      "@      �?       @              �?      �?              �?      �?                       @      d@      &@     �M@       @     �M@      @     �K@      @     �F@       @      D@      �?      &@      �?      &@                      �?      =@              @      �?              �?      @              $@      @      �?       @               @      �?              "@      �?      @               @      �?              �?       @              @       @               @      @                      �?     �Y@      @     �U@              0@      @      (@              @      @               @      @      �?      �?      �?      �?                      �?      @             �j@      B@      ,@      @               @      ,@      @      *@      @      "@      �?       @      �?       @                      �?      @              @       @               @      @              �?       @               @      �?              i@      =@      N@       @      K@              @       @              �?      @      �?      @              �?      �?      �?                      �?     �a@      ;@      �?      @      �?                      @     �a@      8@     �G@      *@      >@      @      >@      @      �?      �?      �?                      �?      =@       @      4@              "@       @      "@      �?      @               @      �?              �?       @                      �?              �?      1@      "@      @      @      @      �?              �?      @                      @      ,@      @      @              @      @      @               @      @      �?      @              @      �?              �?             @W@      &@              �?     @W@      $@      <@             @P@      $@              �?     @P@      "@      O@      @     �F@      @     �F@      @     �D@      @     �B@       @      *@       @      *@      �?       @      �?              �?       @              &@                      �?      8@              @       @               @      @              @       @              �?      @      �?              �?      @                      �?      1@              @       @      @                       @     �@      (@     8�@      (@     0�@      &@     ��@       @     �z@      @     Pu@      @      g@             �c@      @      �?      �?      �?                      �?     �c@       @      @      �?      @                      �?     �b@      �?     �@@      �?      (@      �?      (@                      �?      5@             �]@             �V@      @      G@              F@      @      @       @       @              �?       @               @      �?             �D@       @      4@       @      &@              "@       @      �?      �?              �?      �?               @      �?       @      �?       @                      �?      @              5@             �r@      �?      <@      �?      ;@              �?      �?      �?                      �?     �p@             �S@      @              �?     �S@       @      .@       @              �?      .@      �?       @      �?              �?       @              *@             �O@              �?      �?              �?      �?             �k@             @�@      Z@     �n@     �S@     �n@     �R@      l@     �R@      S@      .@      (@      @      (@      @      "@              @      @       @              �?      @      �?                      @               @      P@      $@     �N@       @     �D@       @     �D@      @      =@      @       @      @      @      @      @      �?      @                      �?              @      @              5@      @      "@              (@      @      @              @      @      @              @      @      �?      @              @      �?               @              (@                      �?      4@              @       @               @      @             �b@     �M@     �U@     �F@      O@      7@      *@      &@      "@      &@       @      @               @       @      @      @      @      @      �?      �?      �?              �?      �?               @                       @      @              �?      @              @      �?      �?              �?      �?              @             �H@      (@      ,@             �A@      (@               @     �A@      $@      &@      @              @      &@      @       @              @      @              @      @              8@      @      ,@      �?              �?      ,@              $@      @      @      @      @      �?              �?      @                       @      @              9@      6@      "@      ,@      �?       @              @      �?      �?      �?                      �?       @      @      @              @      @              @      @      @      @      �?              �?      @                       @      0@       @      0@      @      @              $@      @              @      $@      @      @              @      @      �?      @      �?                      @      @                       @     �N@      ,@      K@      "@      >@      "@              �?      >@       @      1@       @      @              $@       @      "@      @              �?      "@       @      @       @      @      �?      @              �?      �?              �?      �?                      �?      @              �?      @              @      �?              *@              8@              @      @      @              @      @      �?      @      �?                      @       @              5@               @      @       @      �?       @                      �?              @     q@      :@       @      @       @      �?       @                      �?               @     �p@      7@     `d@      6@     �V@      @      4@      @      4@      @      4@       @      @       @      @                       @      0@                      �?              �?     �Q@      �?      ,@      �?      ,@                      �?     �L@              R@      1@      �?      @      �?                      @     �Q@      *@      4@       @      2@      @      "@              "@      @      @      @       @               @      @              @       @      �?       @                      �?      @               @      @              @       @             �I@      @      *@      @      *@       @      @       @      @                       @      $@                      �?      C@       @      6@              0@       @              �?      0@      �?      @      �?              �?      @              *@              [@      �?      2@      �?      2@                      �?     �V@        �t�bub�_sklearn_version��1.2.2�ub.