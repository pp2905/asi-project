����      �!sklearn.neighbors._classification��KNeighborsClassifier���)��}�(�n_neighbors�K�radius�N�	algorithm��auto��	leaf_size�K�metric��	minkowski��metric_params�N�p�K�n_jobs�N�weights��uniform��feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�gender��SeniorCitizen��Partner��
Dependents��tenure��PhoneService��MultipleLines��InternetService��OnlineSecurity��OnlineBackup��DeviceProtection��TechSupport��StreamingTV��StreamingMovies��Contract��PaperlessBilling��PaymentMethod��MonthlyCharges��TotalCharges�et�b�n_features_in_�K�outputs_2d_���classes_�hhK ��h��R�(KK��h�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�_y�hhK ��h��R�(KM:��hB�BЙ                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �t�b�effective_metric_params_�}��effective_metric_��	euclidean��_fit_method��brute��_fit_X�hhK ��h��R�(KM:K��h�f8�����R�(KhCNNNJ����J����K t�b�Bpj       �?                              �?      �?       @      �?                                               @              �?       @fffff�U@fffff�U@      �?              �?             �N@      �?       @      �?       @       @                       @       @              �?       @����̌Z@33333�@      �?                              $@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �3@33333;l@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff3@ffffff3@                      �?      �?      3@              �?                                                                      �?      @������8@�����,{@                      �?      �?      @      �?                       @                                                               @fffff&I@33333#k@                                      �?      �?              �?                                       @       @                       @33333�V@33333�V@      �?                             �P@      �?       @               @       @       @       @                       @                     0Q@���̌_�@                                     �@@      �?       @      �?               @                       @       @              �?       @      Y@33333�@              �?      �?             �F@      �?              �?                       @                       @              �?       @fffff�U@ffff�*�@      �?      �?      �?              P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff�9@333333�@                                      "@      �?       @      �?                                                              �?       @     �R@������@                                      G@      �?       @      �?               @       @                       @      �?      �?       @������W@3333s8�@              �?      �?               @      �?       @      �?               @                                              �?      �?�����)T@fffffʃ@      �?                              7@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333s4@�����~@                      �?      �?     �Q@      �?       @      �?       @               @       @               @       @               @�����Y@3333���@              �?      �?              3@      �?       @      �?                                       @       @              �?       @����̼W@     ��@      �?      �?      �?      �?       @      �?              �?                                       @                      �?      �?�����T@�����;�@      �?              �?              M@      �?       @               @       @       @               @       @       @      �?       @fffff�U@    ��@      �?              �?              R@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����L3@33333c�@                                      "@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?33333s4@�����qb@                      �?      �?      C@      �?                       @       @               @       @       @      �?              �?33333T@����L�@                                      B@      �?              �?                       @       @               @              �?       @33333�U@33333�@      �?                               @      �?              �?                                                              �?       @33333�Q@      b@      �?                              $@      �?                                                               @              �?             `L@     t@      �?                             �O@      �?       @      �?       @       @       @       @       @              �?              �?      Z@����̾�@      �?              �?      �?     �L@      �?              �?               @       @               @       @      �?      �?      �?33333cX@     ޵@      �?      �?      �?      �?     �Q@      �?       @      �?       @       @                       @       @              �?      �?fffffFZ@����|�@                      �?      �?      D@      �?       @      �?                       @       @                              �?       @fffff6U@����Ω@      �?                             �N@      �?       @      �?       @               @               @       @              �?       @����̜Z@ffff&��@                      �?             �@@      �?                               @               @                      �?      �?      �?     �J@33333�@      �?      �?                      @              �?                                                                      �?        3333339@     �Y@              �?      �?              L@      �?       @      �?       @       @       @       @                      �?               @������W@    �_�@              �?      �?              �?      �?       @      �?               @                       @                      �?       @fffff�V@fffff�V@                      �?      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?       @              @������2@������o@      �?              �?      �?      I@      �?       @                               @       @       @              �?      �?       @�����iQ@����L�@      �?                              �?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @�����8@�����8@      �?      �?      �?               @      �?              �?                                                                       @fffff�Q@����̴a@                                      @      �?               @      �?      �?      �?      �?      �?      �?                       @3333334@�����|P@                      �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?       @                     �3@33333�c@      �?      �?                      *@      �?              �?                                       @       @              �?       @     �V@�����Ē@      �?      �?      �?              ;@      �?       @      �?               @       @                       @              �?       @33333�W@fffff��@                      �?      �?     @Q@      �?       @               @                       @                       @              �?33333�N@3333���@                      �?              E@      �?       @      �?                       @       @                              �?      �?�����yU@    �#�@                                      �?      �?       @      �?                                                              �?       @fffff�R@fffff�R@      �?                              0@      �?              �?                                                              �?      �?�����|Q@     ֒@              �?                      �?      �?              �?               @                                              �?       @     @R@     @R@                      �?      �?      4@      �?               @      �?      �?      �?      �?      �?      �?                       @      4@fffffz@                                     �B@      �?              �?               @       @                              �?               @33333T@33333��@                                      @      �?              �?                                       @       @              �?       @fffff�V@�����t|@      �?                              �?      �?              �?                                                              �?       @�����yQ@�����yQ@                                      @@      �?       @      �?                       @               @       @              �?       @fffffVY@������@      �?              �?      �?     �P@      �?              �?               @       @       @       @       @       @                ������Y@    ��@      �?                              I@      �?       @      �?       @       @       @       @       @       @      �?              �?fffff�\@������@      �?              �?              $@      �?       @      �?                                               @              �?       @     PU@fffff��@      �?                              D@      �?                                               @                              �?       @����̌I@�����Y�@      �?              �?              @      �?              �?               @       @                       @              �?       @     �V@     ��@      �?              �?      �?     �I@      �?                       @                       @       @       @      �?      �?        �����S@�������@      �?              �?      �?      E@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     @4@33333��@                      �?      �?      2@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y3@     Ts@              �?                      6@      �?       @      �?                                                              �?        ������R@fffffr�@              �?                       @      �?       @      �?                       @               @       @                       @fffffVY@     d�@                      �?      �?     @Q@              �?               @               @                       @       @      �?      �?������E@33333 �@      �?                              �?      �?                                                                              �?      @fffff&F@fffff&F@      �?                              A@              �?                                                                      �?        �����9@�������@                      �?             �K@      �?              �?       @                               @       @      �?      �?       @     �W@������@              �?      �?              I@      �?       @      �?               @                       @                      �?       @33333V@����Y�@      �?              �?      �?      .@              �?               @                                                      �?        333333>@fffffZ}@      �?              �?      �?      &@      �?       @               @                               @                      �?        �����IP@����̚�@                                     �C@              �?                               @               @       @              �?      �?33333SI@�����ŝ@                      �?      �?      L@      �?       @               @       @                               @      �?                     0Q@�����έ@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?        fffff�3@fffff�3@      �?              �?      �?     �Q@      �?       @               @       @       @       @       @       @       @               @������V@�����@      �?                              :@      �?              �?               @                       @                      �?       @     pU@     Š@              �?      �?              @      �?       @      �?                                                              �?       @fffff�R@������t@      �?              �?      �?      8@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     @4@     |{@      �?                              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     �8@fffffƛ@                                      Q@      �?       @      �?       @       @               @       @       @       @              �?     �[@����Yo�@                      �?      �?     �I@              �?               @                       @                       @                �����A@     ؛@      �?              �?              (@      �?              �?               @                               @              �?      �?33333CU@fffff>�@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @      4@������O@      �?                             �A@              �?                               @               @       @                       @������H@�������@      �?      �?      �?              3@      �?                       @               @               @                                ������P@33333�@                                      A@      �?              �?                                                              �?      �?     �Q@33333�@                      �?               @      �?                       @                       @               @       @              @     `P@����̢�@      �?              �?              C@      �?       @                               @       @               @      �?              �?     @Q@ffff�ڤ@      �?              �?              C@      �?               @      �?      �?      �?      �?      �?      �?       @                ffffff4@     <�@                                     �N@      �?       @               @               @       @       @       @       @              �?����̜U@����L7�@      �?              �?      �?      �?      �?              �?                                       @       @                      @�����IV@�����IV@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff&4@      U@      �?              �?      �?      H@      �?                               @       @                              �?      �?      �?fffff�K@fffff��@      �?              �?              D@      �?       @                       @               @       @              �?              �?     �Q@    �Ӧ@      �?              �?      �?      ?@      �?       @      �?       @               @       @                                       @33333SV@     �@                                     �A@      �?       @      �?                                       @                      �?       @����̜U@33333��@      �?              �?      �?     �A@      �?       @               @       @       @       @                       @      �?      �?�����IQ@����Lt�@                              �?     �P@      �?       @      �?               @               @       @       @       @      �?       @      Z@�����@              �?                      6@      �?                       @               @       @               @              �?      @     pQ@�����%�@      �?                              6@      �?       @      �?                                               @                       @33333�T@33333�@      �?                             �J@      �?       @      �?                                       @                                �����\U@    @��@                                      *@              �?                       @                                              �?       @�����?@     �u@                      �?      �?      6@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     @9@33333[�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      �?����̌4@����̌4@      �?              �?      �?      R@      �?       @      �?               @       @               @       @       @      �?       @������Y@ffff�̼@      �?                              R@      �?       @                       @       @       @       @       @       @      �?        fffff&V@3333�9�@      �?              �?              N@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                fffff&8@�������@      �?              �?      �?      2@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������3@�����du@                              �?      "@      �?                                       @       @       @       @              �?      @�����9R@33333[�@                      �?             �J@      �?              �?                               @       @       @      �?      �?       @�����\W@33333�@      �?                             �M@              �?                                       @       @       @              �?       @������I@�����{�@      �?              �?             �A@      �?       @                       @               @       @              �?      �?       @     @Q@fffff�@                                      *@      �?              �?               @                                      �?      �?      @������R@     2�@                      �?              7@      �?                                       @       @                                       @      K@33333�@                                     �O@      �?       @      �?       @       @       @               @       @                      �?     [@����|�@                      �?      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?      �?              @����̌3@     hr@      �?              �?      �?      =@      �?       @               @                       @       @              �?                33333CQ@����̙�@      �?              �?      �?      6@      �?       @                               @       @       @       @      �?      �?      @������S@     ��@                      �?      �?      R@      �?       @               @       @       @       @               @       @                fffff6T@    ���@      �?              �?      �?     �Q@      �?              �?       @       @       @       @       @               @              �?�����Y@     )�@      �?              �?              @              �?               @       @                                                      @�����A@�����	p@      �?      �?      �?              K@              �?                                                                      �?        33333�8@     S�@              �?                     �J@      �?              �?       @       @               @               @      �?      �?      @     0X@���̌V�@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����L3@fffffb@                                      �?              �?                                                                               @������8@������8@              �?      �?               @      �?              �?                                                              �?       @33333SQ@�����9c@      �?                              @      �?                       @                                       @              �?        33333�M@33333u@                      �?               @              �?                                               @       @                       @�����LF@fffffFX@                                     �O@      �?       @               @       @       @       @       @               @      �?      �?fffff�S@3333s��@              �?                      9@      �?       @      �?               @                               @              �?       @�����lV@�����@                                      <@      �?                       @                       @                      �?              @fffff&K@33333)�@      �?              �?             �M@              �?                                               @       @              �?       @fffff&F@    �դ@                      �?      �?      2@      �?               @      �?      �?      �?      �?      �?      �?                      @33333s4@     Pv@                                      @      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�����L9@�����<]@                      �?              �?      �?               @      �?      �?      �?      �?      �?      �?              �?        �����L4@�����L4@      �?                              @@      �?              �?       @       @       @                       @              �?      �?�����YW@�����F�@                                     �Q@      �?                       @               @       @       @       @       @                fffff�S@3333sյ@      �?                               @      �?              �?                                                                        ����̬Q@33333K�@      �?              �?      �?      :@      �?                                       @                              �?              @�����,I@33333�@              �?                      4@      �?              �?                                               @              �?       @�����\T@fffff�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?fffff�3@������@@      �?              �?      �?      4@      �?                                       @                                      �?       @������H@fffff^�@      �?              �?      �?      E@              �?                       @       @                       @      �?      �?      �?����̌F@�����@      �?              �?      �?      H@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����L:@33333t�@                      �?      �?      N@      �?       @      �?       @       @                       @              �?                ������W@����̳�@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        fffff�4@�����T�@      �?      �?      �?             @Q@      �?       @      �?       @       @                                              �?      �?�����9U@ffff���@      �?                             @P@      �?       @      �?               @       @               @       @       @              �?fffffFZ@������@      �?              �?              3@      �?       @      �?       @       @               @                              �?      �?333333V@fffff!�@      �?      �?      �?             �F@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?33333�8@fffffY�@      �?                              F@      �?                       @                       @       @              �?               @�����YP@������@      �?                               @              �?                                                                              @�����L8@�����9C@              �?                     @Q@      �?       @      �?       @               @       @       @       @       @              �?     �[@���̌+�@                                      C@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@�����1�@      �?                              L@      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @fffff�8@     ؔ@      �?                              $@      �?                                                                              �?       @fffff�F@�����)y@              �?      �?             �Q@      �?       @      �?       @       @       @       @       @       @       @      �?      �?     @\@�����3�@                                     @Q@      �?                       @               @       @       @       @       @      �?      �?����̜T@����L��@      �?              �?      �?      0@      �?                       @       @                                      �?      �?      @������K@fffffΊ@              �?                      *@      �?       @      �?                                               @              �?       @     �T@����̜�@                                       @      �?               @      �?      �?      �?      �?      �?      �?       @              @������4@�����4d@                              �?      2@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����L9@fffffj|@      �?      �?      �?              7@      �?              �?                                       @       @              �?       @����̜V@    ���@      �?              �?      �?     @Q@      �?       @                       @       @       @       @       @       @      �?        �����|T@fffff�@      �?              �?             �P@              �?               @       @               @               @       @      �?        �����yI@fffff��@      �?                              2@      �?       @      �?                                                                      @������R@     ��@              �?      �?              4@      �?              �?                                       @       @      �?      �?             �V@     �@      �?              �?      �?      4@              �?               @               @       @                       @      �?      �?33333�C@33333ˉ@      �?              �?      �?      R@      �?       @      �?                       @                       @       @      �?      �?33333�V@�����o�@                                     �G@      �?       @      �?       @               @               @              �?              �?������W@    @�@      �?                              E@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������3@33333��@                      �?      �?      <@      �?              �?                                               @              �?       @33333CT@33333f�@      �?                              >@      �?              �?       @       @       @                                      �?      �?33333U@33333�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@ffffff4@      �?                              2@      �?              �?                               @                              �?        ������R@33333t�@                      �?              @@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����L3@�������@                                      6@      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@33333c}@      �?                               @      �?              �?                                                                      �?����̬Q@fffff�a@      �?                              @      �?                               @               @       @                      �?             �O@fffffFl@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@fffff��@      �?              �?      �?      R@      �?       @               @       @       @       @       @               @      �?        fffff6T@3333s_�@      �?      �?      �?              $@      �?       @      �?                                               @              �?       @������U@33333Ŋ@      �?              �?      �?     @Q@      �?       @               @               @       @       @       @       @                ������U@����2�@      �?                      �?      $@      �?       @       @      �?      �?      �?      �?      �?      �?                      �?������8@������k@      �?                      �?      ?@      �?       @                       @               @       @       @      �?      �?      @������S@fffff7�@                                      @      �?              �?                                                                       @������Q@     �q@      �?                              �?      �?                                                       @                      �?      @     �J@     �J@      �?              �?              (@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������3@     Hi@      �?                              R@      �?       @      �?               @       @               @       @      �?      �?       @�����<Z@����Lx�@      �?      �?                      6@      �?       @      �?                               @       @                      �?             �V@fffffڝ@                                      4@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �3@fffff2y@      �?                             �I@      �?       @      �?               @       @       @                              �?       @fffff�U@     y�@                                      2@      �?       @      �?                               @       @                      �?       @fffffV@33333��@      �?      �?      �?      �?     �P@      �?       @      �?               @       @       @       @       @      �?      �?       @�����[@����Y��@      �?              �?      �?      E@      �?       @               @       @                       @                      �?        �����YQ@������@                                       @      �?               @      �?      �?      �?      �?      �?      �?       @              @      4@33333�a@      �?                              C@      �?       @      �?                       @       @       @              �?                     �W@33333+�@                                      �?      �?              �?                                                              �?       @�����LQ@�����LQ@      �?              �?             �J@              �?                       @       @       @       @       @      �?      �?       @�����9N@    ��@                      �?             �O@      �?              �?       @               @                              �?      �?      �?�����IT@    �h�@      �?              �?      �?      @      �?                       @                                              �?      �?       @     �H@����̴t@                              �?      .@      �?              �?                                                                             @Q@fffff�@      �?                             �I@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �8@fffffJ�@              �?      �?              *@              �?                                               @       @                       @fffff�F@�������@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@     �3@                                      O@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?3333333@�������@                      �?             �A@      �?                               @               @                                       @�����lL@fffff�@                                      �?      �?              �?               @                       @                               @33333U@33333U@                      �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�3@33333��@      �?              �?      �?      *@      �?                                                                                        ffffffF@�����y�@                      �?              5@      �?              �?                       @       @                      �?               @������S@�����9�@      �?                      �?      J@      �?       @               @       @               @       @       @       @      �?      @�����IU@�����m�@      �?              �?      �?     �E@      �?                       @               @       @       @       @       @      �?      �?������S@33333ݫ@      �?                               @              �?                       @       @       @                              �?      �?333333D@�����IS@      �?                              0@      �?       @      �?               @                                              �?      @33333#T@�������@      �?              �?              L@      �?       @      �?               @                       @       @      �?              �?33333Y@3333s�@      �?              �?      �?      N@      �?               @      �?      �?      �?      �?      �?      �?       @              @����̌4@33333Ԓ@      �?      �?      �?              8@      �?       @      �?       @                                                      �?       @fffff�S@     ��@                                      $@      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�4@     �n@      �?              �?              7@      �?                       @                                       @              �?        ������M@     ��@      �?                              O@      �?       @      �?       @       @               @               @      �?               @     �Y@    @��@                      �?      �?     �M@      �?       @               @       @               @                      �?              @     `P@�������@      �?                              2@      �?               @      �?      �?      �?      �?      �?      �?                      @     @3@������t@      �?              �?      �?     @P@      �?       @      �?       @       @       @       @                       @              �?33333�W@    ���@      �?                               @      �?              �?                                                                      @����̬Q@fffff&`@      �?              �?             �H@      �?       @      �?       @       @                       @                      �?        fffffvW@����}�@      �?      �?      �?              C@      �?       @      �?               @       @               @       @              �?       @fffff�Y@fffffR�@      �?                              �?              �?               @                                                              @33333�=@33333�=@                      �?             �Q@      �?       @      �?       @       @                       @              �?              @������W@3333�Ⱥ@                              �?      @      �?       @      �?               @                       @                              @ffffffV@fffff�v@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@����̌;@      �?              �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?        33333]@    �4�@      �?                              >@      �?       @      �?                               @               @              �?      �?�����yV@����LF�@      �?              �?      �?     �A@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@fffffz�@      �?              �?              N@      �?       @      �?               @       @               @                      �?       @     �W@ffff�n�@                              �?      A@      �?       @      �?       @       @       @       @       @       @       @      �?      �?�����	]@�����ծ@                      �?             �H@      �?               @      �?      �?      �?      �?      �?      �?      �?                33333s4@33333'�@      �?                      �?      1@      �?                               @       @       @       @       @      �?               @fffff6T@����̗�@      �?                              "@              �?               @               @       @               @      �?              @ffffffI@������|@                      �?      �?      :@      �?              �?       @       @                                                       @�����|T@����,�@      �?      �?                      J@      �?       @      �?                                                              �?        �����<R@    ��@      �?              �?             �I@      �?       @      �?       @               @       @       @       @      �?      �?       @33333�[@����YX�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @����̌3@����̌3@      �?              �?      �?      �?      �?              �?                                       @       @              �?       @fffff�V@fffff�V@                                      =@      �?               @      �?      �?      �?      �?      �?      �?       @              @ffffff3@     R�@      �?              �?             �M@      �?       @      �?       @       @       @               @       @      �?      �?       @������[@����0�@      �?      �?                      5@      �?       @      �?               @       @               @       @              �?       @fffffZ@3333���@                                      *@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @ffffff4@�����Tp@                                     �A@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����5@     (�@                                      �?      �?       @      �?                                               @              �?      @�����\U@�����\U@                                      H@              �?               @       @                       @                      �?       @ffffffF@����q�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@33333M@                                      @      �?       @      �?               @                                                        �����|S@�����s@      �?                              5@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�����Y4@33333kz@      �?              �?      �?     �P@      �?       @               @               @               @       @       @      �?       @������S@fffff��@                      �?             �N@      �?       @      �?               @                       @       @       @      �?        33333CY@    @S�@      �?                              P@      �?       @                       @       @       @       @       @       @              �?33333�U@���̌ �@      �?              �?      �?      "@      �?              �?               @               @       @       @              �?       @     `Y@�����V�@              �?      �?             @P@      �?       @      �?       @               @               @       @                             PZ@fffff��@      �?              �?             �B@      �?       @               @               @               @       @      �?              @     �S@�������@                      �?      �?     �A@              �?                                       @       @              �?              @33333sD@fffff��@      �?      �?                      �?      �?       @      �?                       @               @                      �?       @333333V@333333V@      �?              �?              ,@      �?                               @       @       @       @       @       @              @�����|T@     w�@      �?              �?      �?      R@              �?               @       @       @       @       @       @       @      �?      �?333333P@    �o�@              �?                       @      �?       @      �?                       @                                      �?       @33333�S@������b@              �?                      @      �?              �?               @                       @                      �?       @�����,U@     �x@      �?                              6@      �?       @      �?       @                               @       @              �?       @     0Y@     ^�@      �?              �?              >@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@33333�@      �?              �?      �?     �G@      �?       @      �?               @                       @       @              �?       @fffff�X@ffff&��@                      �?              9@      �?              �?                       @                                      �?       @fffff�R@     �@      �?                              �?      �?                       @                                                      �?      @     `I@     `I@      �?              �?      �?     �I@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @33333�8@     �@                              �?      :@      �?       @                                                                      �?      @     �H@�����Ɠ@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����4@      �?                              K@      �?       @      �?               @                                              �?        fffff�S@    @԰@                      �?             �M@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����Y4@     ̓@                      �?      �?     �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�����8@fffff>�@      �?                      �?      @      �?       @      �?                       @                       @                       @fffff�V@�����p@              �?                      @      �?              �?                                                              �?      @33333CQ@     �s@      �?              �?      �?      =@      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�4@�����v�@                                      @      �?                       @       @                                                      @33333�K@fffff.t@                                     �J@      �?              �?               @       @       @               @      �?      �?      �?����̜W@    ���@      �?                              R@      �?       @               @       @       @       @       @       @       @                      W@    ��@                      �?      �?     �@@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @     �8@fffff"�@      �?      �?      �?             �@@      �?       @      �?                                       @       @              �?       @     �W@����C�@      �?                             @Q@      �?       @               @       @       @       @               @      �?      �?      �?fffff�S@3333s�@      �?                              �?              �?                                               @       @              �?      @fffff�F@fffff�F@      �?              �?      �?     @Q@      �?       @      �?               @       @               @       @       @      �?       @     @Z@    ���@      �?                              "@      �?                                                                              �?      @333333F@fffff�u@                                      @      �?              �?                                               @              �?       @������S@     �s@                                     �Q@              �?               @               @       @       @       @       @      �?        �����,M@    @v�@                              �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @     �3@     |�@      �?              �?      �?      7@      �?                       @                       @                      �?              �?������L@fffff=�@                      �?      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@�����
�@      �?              �?              ;@      �?                       @                                              �?              �?�����YH@     7�@      �?                              A@      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@������@      �?      �?      �?             �P@      �?                       @       @               @                      �?      �?        �����yN@fffff�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                       @     @3@33333\@                                      @      �?                                                               @              �?       @     �K@fffffFu@                      �?      �?      0@      �?              �?               @       @               @                      �?      �?�����\V@     Y�@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @3333334@fffff�X@              �?      �?             �Q@      �?       @               @       @       @       @               @       @      �?        ����̬T@33333Ƕ@                                     �P@      �?       @      �?       @       @       @       @               @              �?        fffff�Y@     ù@              �?      �?             �K@      �?              �?                       @       @       @               @              �?333333V@����LŲ@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff6]@����َ�@      �?                              G@      �?               @      �?      �?      �?      �?      �?      �?       @                �����4@     0�@                      �?              P@      �?              �?       @               @               @       @       @      �?             �X@������@                      �?              ,@      �?              �?       @       @               @       @       @      �?              @�����|Z@������@      �?      �?                      &@      �?       @      �?               @       @       @       @       @              �?       @������[@33333|�@      �?      �?      �?             �E@      �?       @      �?               @                       @       @              �?       @     @Y@fffff$�@                                       @      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333s4@�����9E@      �?              �?      �?       @      �?                                       @                                      �?       @fffff�I@������y@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @ffffff3@�����e@      �?                              "@      �?                       @               @       @               @              �?             Q@������@      �?                      �?     �C@              �?               @                       @       @              �?                fffff�F@fffff��@                              �?      7@      �?                                               @                      �?      �?       @������H@fffff}�@                      �?              �?      �?              �?                                                              �?      @�����YQ@�����YQ@      �?      �?      �?              &@      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@     �j@      �?                              5@      �?       @      �?                                                              �?       @�����lR@�����Z�@                                     @P@      �?       @      �?               @               @       @       @      �?      �?        33333CZ@    @X�@      �?                             �P@      �?                                               @                       @                fffffFI@33333x�@      �?              �?              L@      �?              �?                                       @       @                      @�����lV@3333�X�@              �?                      @      �?       @      �?                                       @       @              �?       @33333�W@33333�z@      �?      �?      �?              F@              �?                       @                                              �?       @�����Y>@�����>�@      �?              �?              R@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�3@�����7�@                      �?             �G@      �?       @      �?                       @               @       @              �?       @      Y@����c�@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?�����I]@    ���@      �?                              �?      �?                       @                       @                              �?       @������J@������J@      �?              �?              L@      �?              �?                                               @      �?      �?       @�����9T@    �ͱ@      �?              �?      �?      0@      �?               @      �?      �?      �?      �?      �?      �?                       @fffff&4@�����Uu@      �?              �?              E@      �?       @      �?                       @       @       @       @              �?        ������Z@3333���@      �?                      �?     �Q@      �?       @      �?       @       @                                      �?      �?      �?�����\U@3333�@                                      G@      �?              �?               @       @       @       @       @       @      �?        �����Z@33333(�@      �?                              H@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@     ��@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�4@     �L@                      �?              <@      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@fffff��@      �?              �?              R@              �?               @       @       @       @       @       @       @      �?       @�����,P@������@              �?                     �D@      �?              �?                       @       @       @       @      �?      �?        fffffFY@fffff`�@              �?      �?              8@      �?       @      �?                                       @       @              �?       @33333cW@������@      �?      �?      �?              *@      �?              �?               @       @               @       @              �?       @     �X@fffffW�@                      �?      �?     �K@      �?       @      �?       @                               @       @      �?              @�����9Y@�����H�@      �?              �?              >@      �?       @                                                                               @33333�H@����̇�@                      �?              G@      �?       @               @                                                                     �K@ffff�S�@      �?      �?                      7@      �?       @      �?               @       @               @       @              �?       @������Z@     g�@                                      @      �?              �?                       @               @       @              �?       @fffff�W@33333��@      �?      �?                     �P@      �?       @      �?                       @               @       @              �?      �?�����YY@������@                      �?      �?      $@      �?                                       @       @                                      �?������K@����̂�@                                      :@      �?       @      �?                       @                                      �?       @�����,T@     "�@      �?      �?      �?              @      �?       @      �?                                                              �?       @������R@fffff��@                                      @      �?                                               @       @       @              �?      �?     �Q@�����,|@                                      Q@              �?                       @               @               @                       @�����yF@3333��@                      �?              .@      �?              �?                                       @       @                       @�����	V@fffff��@                      �?      �?      @      �?       @                       @               @                              �?      @     @M@33333l@      �?                              7@      �?       @      �?                               @       @                      �?       @fffff�V@�����\�@      �?              �?      �?      9@      �?              �?                                       @       @      �?      �?       @������V@33333�@      �?                              "@      �?       @      �?                                                              �?       @fffff�R@33333��@              �?                      4@      �?       @                                                       @              �?      @������N@fffffY�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?       @3333334@������K@              �?      �?              1@      �?       @      �?                                       @       @              �?       @33333#W@�����:�@      �?                             �@@      �?              �?               @               @                       @                fffff&T@33333��@                      �?             �B@      �?       @      �?       @               @       @               @      �?      �?       @������X@33333U�@      �?                              �?      �?                                                                              �?       @     `F@     `F@                              �?      3@      �?       @               @       @               @       @                      �?      @������R@fffff~�@              �?                     �C@      �?       @      �?                       @               @       @              �?       @     �X@     ��@      �?              �?             �G@      �?       @       @      �?      �?      �?      �?      �?      �?                       @ffffff9@�����̑@                                      @      �?                                               @                              �?        ffffffI@����� r@      �?              �?      �?     �N@      �?       @      �?       @       @                       @       @      �?      �?       @     �Z@3333���@                                      =@              �?                       @                                              �?       @������>@�����@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?                      @      4@33333;q@                      �?              1@      �?       @      �?                                       @       @                       @fffff&W@����̮�@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�4@     �b@      �?              �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @ffffff9@�������@      �?                              C@      �?       @      �?       @       @                       @       @      �?      �?       @fffff6Z@    �^�@      �?                             �P@      �?       @      �?               @                               @                      �?�����YV@ffff�X�@                      �?              $@      �?               @      �?      �?      �?      �?      �?      �?              �?      @����̌4@     �o@      �?              �?      �?       @      �?              �?                                       @       @              �?        33333cV@�����1g@                      �?      �?     �A@      �?                       @                       @                      �?      �?        �����yK@     �@                      �?              L@      �?              �?       @       @       @               @       @      �?      �?      �?ffffffZ@ffff���@              �?      �?              .@      �?       @      �?                       @       @                              �?       @33333�T@33333��@                      �?              Q@              �?               @               @               @       @      �?      �?       @333333K@����L�@              �?      �?             �Q@      �?       @      �?       @       @       @       @                       @      �?      �?fffffX@3333�n�@      �?                              5@      �?                       @               @               @                                fffffVP@�����A�@      �?              �?      �?     �P@      �?       @      �?       @       @       @               @       @      �?      �?       @33333�[@����:�@              �?      �?              I@      �?       @      �?               @       @               @                      �?       @33333�W@3333��@              �?                      @              �?                                                                               @�����L9@     pS@                      �?      �?      @      �?                               @               @                                      @     @L@33333cm@      �?                              .@      �?       @      �?                                       @       @              �?       @fffffVW@�������@      �?              �?              R@      �?       @      �?               @       @       @       @       @       @      �?       @�����[@�������@      �?                              G@      �?               @      �?      �?      �?      �?      �?      �?       @               @33333�3@fffffX�@              �?                       @      �?       @      �?                                                              �?       @     �R@     �@                                      @@      �?       @      �?               @       @               @       @      �?      �?      �?33333Z@3333���@      �?      �?                      8@      �?       @      �?               @                       @       @              �?       @     PY@����L�@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?       @                33333�3@     �@                                      @      �?              �?               @                       @       @                       @������W@fffffRr@                      �?      �?     �Q@      �?                       @       @       @       @                       @              �?33333P@ffff挱@      �?              �?             �P@      �?                       @       @               @               @       @      �?      �?�����LQ@ffff�?�@      �?              �?      �?      &@      �?              �?                                       @       @                       @fffff�V@������@              �?                      @      �?              �?                       @               @                      �?       @fffff�U@fffff�k@      �?                               @      �?              �?                                                              �?      @fffff�Q@�����:�@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        33333�\@    @��@      �?                               @      �?                       @                                                      �?       @fffff�G@�����W@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@      M@                                     �P@      �?                       @       @       @                               @      �?        33333�N@ffff�b�@      �?              �?      �?      ,@      �?                       @       @                               @       @      �?        33333�N@fffff|�@                                      (@              �?                       @       @       @       @       @      �?               @33333SN@fffff:�@      �?              �?              @              �?                       @                       @       @              �?       @fffffFH@      i@              �?                      R@      �?       @      �?       @       @       @       @               @       @      �?        ������Z@    �D�@      �?      �?                     �Q@              �?               @       @                       @       @      �?      �?       @�����9L@3333�"�@                      �?             @P@      �?                       @       @       @                       @       @                     �Q@33333"�@      �?                              9@      �?              �?                                                                       @     pQ@fffff�@                      �?             �I@      �?                       @       @               @                      �?      �?             @N@����L��@              �?      �?             �P@      �?       @                       @       @               @              �?      �?        fffff�Q@����ق�@                      �?      �?     �@@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?fffff&8@fffff�@      �?                              8@      �?                                       @                                      �?      @������H@33333?�@      �?      �?                      K@      �?                                       @       @               @      �?                     PP@ffff擫@      �?              �?      �?      *@      �?                                                       @       @      �?      �?       @     0P@�����j�@                      �?      �?      M@      �?              �?               @       @               @                      �?       @33333�V@ffff���@                      �?             �H@      �?       @               @       @       @                       @      �?               @33333�Q@���� �@                      �?              :@      �?       @               @       @       @       @       @       @      �?      �?      �?fffff�V@�����@                      �?             �F@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �9@33333��@                      �?             @P@      �?       @      �?       @       @               @       @              �?      �?        �����	Y@    ��@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@�����\W@      �?                              @              �?                                                                               @     �8@����̼P@      �?                             �C@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@33333��@              �?                      F@      �?              �?               @       @                       @      �?              �?�����IV@    �-�@                      �?              "@      �?              �?                       @                                      �?             �R@33333�@      �?              �?      �?      B@      �?                       @       @                                      �?              @33333�J@fffffM�@      �?              �?              @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y3@33333�_@                                      .@      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@33333t@              �?                     @P@              �?                       @       @               @       @       @      �?             �J@�����{�@                      �?             �Q@      �?       @               @       @       @       @       @       @       @               @fffff�V@ffff榸@      �?              �?      �?     �Q@      �?       @               @       @       @       @       @       @       @              �?�����yV@ffff&9�@      �?              �?      �?     �Q@      �?       @               @       @       @       @       @       @       @      �?      @     �V@�������@                      �?      �?      �?              �?               @                                                                     �>@     �>@                                      (@      �?                                                                              �?       @fffff�F@�����X�@                      �?               @      �?                                                                              �?      �?�����LF@33333#T@                                      @      �?              �?                                       @                      �?       @     �S@fffff�r@                      �?      �?     �F@      �?       @      �?       @       @                       @       @              �?       @�����IZ@ffff�z�@                      �?              R@      �?       @      �?       @       @       @               @               @                �����)Y@������@      �?                              A@      �?       @      �?       @       @       @       @       @       @      �?              �?     ]@����v�@      �?              �?              E@      �?       @      �?       @               @                       @              �?       @������W@33333]�@                                      =@              �?                                       @                              �?       @333333?@������@      �?      �?      �?              @      �?       @      �?                                       @       @              �?       @fffff�W@�����xq@      �?                              ?@      �?              �?                       @       @       @       @       @                ������X@�����K�@      �?                              �?      �?                                                               @              �?       @     �K@     �K@              �?      �?              O@      �?       @      �?               @       @               @              �?      �?      �?�����|X@���̌0�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @      4@      4@                                      1@      �?       @                               @       @       @                      �?      @     @Q@     P�@      �?                              @@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����4@�����3�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����L4@�����L4@      �?              �?      �?      <@      �?       @      �?       @       @                       @       @      �?               @fffff�Z@�����>�@                                      �?      �?       @      �?               @                                              �?      @������S@������S@                      �?      �?      H@      �?              �?       @               @               @       @      �?      �?        ������X@33333q�@              �?      �?             @Q@      �?       @      �?               @               @       @       @       @              �?�����YZ@3333�V�@              �?                      E@      �?       @                               @                                               @33333�K@    ��@                                      �?              �?                                                                      �?      @�����9@�����9@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@fffff�C@              �?      �?              :@      �?              �?               @                               @                       @�����<U@    ��@                      �?      �?      ;@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@�����0�@                      �?      �?     �E@      �?       @      �?                       @                       @              �?        33333#W@     ��@      �?                              �?      �?              �?                                       @                      �?       @33333�S@33333�S@              �?                      �?      �?              �?               @                               @              �?       @     �U@     �U@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@fffffS@      �?                              �?      �?                               @                                              �?      @33333I@33333I@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff&4@fffff&4@                      �?      �?      R@              �?               @       @       @       @       @       @       @                �����P@     ��@                                      @      �?                                                                              �?      @fffff�F@fffff�h@              �?      �?      �?      R@      �?       @               @       @       @       @       @       @       @              �?�����W@    @(�@                                      �?      �?              �?                                                              �?       @fffff�Q@fffff�Q@      �?              �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @              �?     �\@����L��@              �?                      3@      �?              �?       @       @               @       @       @              �?      @     @Z@     ]�@                      �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?      �?               @������3@�����d@      �?      �?      �?              �?              �?                                                                               @�����9@�����9@      �?      �?                     �O@      �?       @      �?       @       @       @               @       @              �?        �����Y[@3333sw�@      �?                              :@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@����̔|@      �?              �?      �?     �P@              �?                                       @       @       @       @                fffffFI@����I�@      �?                              6@      �?                       @                       @                                      @����̌K@�������@                                      K@              �?               @                       @               @      �?                �����F@fffff��@      �?              �?              N@      �?                       @       @               @                       @      �?      @����̬N@fffffl�@                              �?      @      �?               @      �?      �?      �?      �?      �?      �?              �?        �����4@     `U@                                      �?      �?                                                                              �?      @      F@      F@      �?                             �P@              �?               @               @       @       @              �?      �?        ����̬H@3333��@              �?                      I@      �?       @      �?       @       @                                              �?       @������T@3333��@      �?                              (@      �?              �?                                               @              �?        ������S@�����M�@      �?              �?      �?     �@@      �?                       @               @               @       @      �?              �?     �R@�����*�@              �?                      =@      �?       @      �?                               @       @       @                       @������X@    �]�@      �?                              @              �?                                               @       @              �?       @fffffFF@������e@      �?                      �?      D@              �?               @       @               @                      �?              @      D@33333p�@      �?                             �I@      �?              �?       @                               @              �?              @fffff�U@ffff&��@                      �?      �?      *@      �?                                                               @                       @������K@������@      �?      �?      �?             �Q@      �?       @      �?       @       @       @               @       @              �?       @     �Z@���̌!�@                      �?             �P@      �?       @               @       @       @                               @                ������P@    @�@              �?      �?              I@      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @3333339@33333i�@                                     �D@      �?       @      �?       @       @       @       @       @       @              �?             �\@3333s��@                      �?      �?      @      �?                       @       @       @               @              �?               @�����\Q@������}@                                      ,@      �?              �?                       @                                               @fffff�R@������@      �?                              Q@      �?       @      �?               @       @       @       @       @      �?               @�����[@���̌�@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@33333�b@                                      @              �?               @       @                                              �?       @33333�@@33333;a@      �?      �?      �?             �A@      �?       @      �?                       @                              �?      �?        ffffffT@    ���@              �?                      A@              �?                       @       @               @       @              �?       @      L@����̗�@                                      @      �?              �?               @                       @                      �?      @33333SU@33333Gz@                                     �G@      �?       @      �?               @       @               @       @              �?       @������Z@3333��@                                      5@      �?                       @       @               @       @               @              �?33333�Q@fffffӗ@      �?                              �?      �?                                                                              �?      @33333sF@33333sF@                      �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�4@33333)�@      �?                             �A@      �?       @      �?       @               @       @       @       @       @      �?       @�����<[@     s�@      �?              �?      �?      *@      �?              �?       @                                       @                       @33333U@33333�@      �?                              ?@      �?              �?               @                       @       @              �?       @     �W@fffffF�@      �?                              ?@      �?              �?               @               @                              �?       @����̜S@����L�@      �?                              @      �?       @      �?               @       @               @       @                      @������Z@������s@      �?                              3@      �?       @      �?       @               @                                      �?       @     0U@�����ϙ@                                      �?      �?              �?                                                              �?       @fffff�Q@fffff�Q@              �?      �?              E@      �?       @      �?       @               @               @       @      �?      �?        �����LZ@ffff&��@      �?                              R@      �?       @      �?               @       @       @       @       @       @                �����L[@����Lƾ@      �?              �?      �?      N@      �?                       @       @       @       @                      �?      �?        fffffvP@�������@                                      �?      �?              �?               @       @                                      �?       @33333�T@33333�T@                      �?      �?      B@      �?               @      �?      �?      �?      �?      �?      �?       @                     @4@�����o�@      �?              �?      �?     �E@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     @8@�����א@                      �?      �?      "@      �?       @                       @                                              �?      @fffff�K@33333S@                      �?              ;@      �?              �?       @                       @       @       @      �?      �?      �?�����yY@����L�@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������8@fffff?�@      �?                             �A@      �?       @      �?                                       @                               @������T@ffff�@�@      �?      �?      �?              A@      �?              �?                                                                      �?33333�Q@3333���@                      �?             �L@      �?                       @       @               @       @               @      �?      �?fffff�Q@ffff��@                      �?      �?     �H@      �?       @      �?               @                       @       @      �?              @�����Y@�����M�@                                      (@      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@33333�k@      �?                              R@              �?               @               @       @       @       @       @      �?      �?������N@    @&�@      �?              �?      �?     @P@      �?       @               @       @       @                       @      �?              �?�����R@�����-�@      �?              �?      �?      ;@      �?       @      �?       @       @               @       @                               @     0Y@����ӥ@      �?              �?              @      �?              �?                                       @                      �?       @fffffT@fffff6s@                      �?              R@      �?       @      �?               @       @               @       @      �?      �?       @fffffVY@ffff&��@      �?              �?              R@      �?       @      �?               @       @       @       @       @       @      �?      �?fffff�[@33333�@      �?              �?              5@      �?       @      �?                       @       @       @       @              �?       @fffff�Z@ffff擡@      �?              �?      �?      M@      �?       @      �?                       @       @               @       @                fffff�W@ffff���@      �?              �?             �@@      �?                                                                              �?      �?fffffFF@fffffږ@                      �?              *@      �?                                                                      �?               @fffff�E@33333��@                                      �?      �?              �?                                               @              �?       @�����|T@�����|T@                      �?      �?     �N@      �?       @               @       @       @       @               @      �?      �?       @������S@���̌Բ@      �?                              &@      �?                                                                                      �?������F@     �~@              �?                      C@      �?                       @       @                                              �?      �?33333�L@����L��@                      �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @                33333�3@�����ӕ@      �?                              >@      �?                       @       @               @       @              �?               @������Q@     �@      �?                              9@      �?              �?                       @       @       @       @       @                33333�X@     ��@                                      *@              �?                               @               @       @                       @33333�H@33333K�@      �?                              E@      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�����9@����̮�@                                      "@      �?              �?                       @                       @              �?      �?33333SU@33333k�@      �?              �?              *@      �?       @      �?                       @               @       @              �?      �?     �Y@     <�@                      �?             �O@      �?       @      �?               @       @       @       @       @              �?       @     0[@3333�׺@      �?              �?      �?      C@      �?       @      �?                       @               @       @              �?      �?�����IY@fffff�@      �?              �?      �?      A@              �?               @                                              �?                ffffff>@33333U�@      �?                              .@      �?              �?                       @       @       @       @              �?       @fffffVY@�����G�@                      �?              R@      �?       @               @       @       @       @       @       @       @                      W@fffffJ�@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?        33333�\@3333st�@      �?              �?      �?      G@      �?                       @               @       @       @       @       @              @     @T@3333��@      �?              �?      �?      R@      �?              �?       @       @       @       @       @       @       @                ������[@����a�@                                      �?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @     �9@     �9@      �?              �?             �Q@      �?       @               @       @               @                       @                �����IP@    �I�@                              �?      9@      �?               @      �?      �?      �?      �?      �?      �?                      �?�����4@33333{}@              �?                     �E@      �?              �?       @       @               @       @       @              �?      �?�����	[@3333���@      �?              �?      �?      &@      �?              �?                                       @                      �?             �S@     $�@      �?              �?      �?      R@              �?               @       @       @       @       @       @       @      �?      �?     PP@�����~�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      �?�����L4@�����L4@      �?                              �?      �?              �?                                                              �?       @fffffvQ@fffffvQ@      �?              �?      �?      @      �?                               @       @                                      �?      @fffff�K@     Dt@      �?                              R@      �?       @               @               @       @       @       @       @              �?33333U@����m�@                      �?      �?      H@              �?                                       @                              �?      �?     �=@33333<�@      �?              �?      �?     �J@      �?                       @       @               @       @               @      �?      @�����lQ@33333#�@                                      @      �?              �?       @               @       @               @              �?        ������W@333333x@                      �?              @      �?              �?                                                                       @�����|Q@fffff�t@                      �?              8@      �?              �?               @       @               @       @              �?      �?33333�X@3333���@                                       @      �?                               @               @       @                      �?       @�����\P@�����S�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@     �3@                      �?      �?      M@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff&9@�������@                              �?     �D@      �?       @      �?               @                       @                      �?              V@����z�@      �?                      �?      L@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @������8@�����@�@      �?              �?              R@      �?       @                       @       @       @       @       @       @      �?        �����IU@33333��@                      �?               @      �?              �?                                                              �?      �?������Q@�����Yc@      �?              �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @�����Y4@     >�@      �?              �?              7@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����L3@33333c~@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@      �?                              9@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?             �3@fffff"�@      �?                              @      �?              �?               @                       @                      �?       @fffffVU@33333�~@      �?                             �B@      �?       @               @       @       @       @                      �?               @������P@������@      �?              �?      �?     @Q@      �?       @      �?                               @       @       @       @      �?       @fffff�X@3333sȺ@      �?                              0@              �?               @       @       @       @       @               @              @�����lK@33333��@      �?                               @      �?       @      �?                                               @                              U@33333��@                                      E@      �?               @      �?      �?      �?      �?      �?      �?       @      �?             �4@�����c�@      �?      �?                      @      �?                                                                                      �?�����YF@     Hq@                                      @      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�3@fffff6]@      �?      �?                     �G@      �?       @      �?                                       @                      �?      �?33333�U@333333�@      �?      �?                      ?@      �?       @      �?               @                       @                      �?       @����̬V@����L:�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@�����4@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @                33333s3@     ^�@                      �?              B@      �?       @      �?       @       @       @       @               @       @      �?      �?33333�Z@�������@                                     �P@      �?       @      �?       @       @       @               @                      �?      �?����̼Y@    @�@                      �?              E@      �?       @               @       @               @                              �?      �?������P@�����O�@                      �?              0@      �?       @      �?       @       @       @                                               @����̬V@�����{�@              �?      �?              H@      �?       @      �?       @       @       @       @       @       @                       @�����\]@ffff�>�@                                      *@      �?                       @                       @                      �?              @33333�K@333337�@      �?                              >@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@fffff��@                                     �G@      �?                                       @       @       @       @       @              @����̜R@�����l�@      �?      �?      �?              F@      �?       @      �?               @                               @      �?              @�����V@����̑�@                      �?             �H@              �?                       @               @       @       @      �?      �?      �?fffff&L@33333��@                                      2@              �?               @       @               @                      �?      �?      @�����D@�����?�@                              �?      ,@      �?       @      �?       @                       @                              �?      @     �U@333330�@      �?              �?      �?      R@              �?               @       @       @                               @              �?     @C@     ��@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?       @                33333�3@33333��@                      �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333�8@33333J�@      �?      �?      �?              K@      �?       @      �?                                                                             �R@����L��@      �?                              @      �?       @      �?                                                              �?       @fffff�R@������p@              �?      �?              N@      �?              �?       @       @       @       @       @       @       @      �?             �[@����Y�@                      �?              J@      �?                       @               @               @              �?      �?      @33333P@33333��@      �?                              J@      �?              �?               @       @       @       @       @      �?      �?             @Z@�����2�@      �?              �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @               @����̌4@33333b�@      �?      �?      �?      �?      R@              �?               @       @       @       @       @       @       @      �?        333333P@����Y|�@                                      .@      �?                       @       @       @       @       @       @                      @�����U@fffff�@      �?                             �K@      �?       @                               @               @       @       @      �?        33333sS@����Y�@      �?                              J@      �?              �?       @               @               @              �?               @     �V@����L��@      �?                              I@      �?              �?       @       @       @       @                      �?      �?      �?fffff�V@3333sű@                                      .@      �?                                                       @              �?              @33333L@33333�@      �?                              2@      �?       @               @               @               @                              @     `Q@�������@      �?                      �?      *@      �?              �?                                       @                      �?      �?33333�S@�����'�@      �?              �?              J@      �?       @      �?               @               @               @              �?      �?������W@fffff�@                                      O@      �?       @                       @       @       @       @       @       @                      U@33333I�@      �?                             �C@              �?               @       @               @       @                      �?      �?�����yH@fffffc�@      �?              �?              (@      �?              �?       @       @       @                                      �?       @fffff&U@33333��@      �?                              O@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�����4@�����ƒ@                                      6@      �?       @      �?                                                      �?      �?      �?      S@fffffޛ@                                      �?      �?              �?                                                                       @     �Q@     �Q@              �?                      R@      �?       @      �?               @       @       @       @       @       @      �?        fffff[@����^�@      �?              �?      �?      6@      �?                                               @                              �?       @����̌I@�����C�@                                      F@      �?              �?               @       @               @                      �?      �?�����	V@fffff
�@      �?      �?      �?             �H@      �?       @      �?               @                               @                      �?33333�V@    @ñ@      �?              �?      �?      O@      �?                       @               @       @               @      �?              �?������Q@����L��@              �?                      2@      �?                               @                                              �?      �?������H@     �@                      �?      �?     �D@      �?              �?                       @               @       @              �?        ������W@     �@      �?                              �?      �?              �?                                                              �?       @fffffVQ@fffffVQ@      �?                              �?      �?                                       @       @                                      @fffff�K@fffff�K@      �?                              R@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������4@�����ė@      �?              �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@fffff�t@      �?                             �P@      �?                       @               @                       @       @                33333cP@���̌	�@                                      8@      �?       @      �?               @       @               @       @              �?       @�����	Z@����L}�@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?                             �3@�����Ib@                      �?              R@      �?       @      �?       @       @       @       @                       @      �?             @X@33333��@      �?              �?      �?      8@      �?       @               @                       @       @       @                             @T@fffff�@      �?                             �B@      �?       @               @       @       @       @       @       @      �?      �?        fffff�V@����L=�@                      �?      �?      <@      �?              �?       @                                       @      �?      �?        fffff�T@�����!�@                      �?      �?     @Q@      �?                               @       @       @                      �?                ����̌M@3333�&�@                      �?      �?      N@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?     @3@     =�@      �?      �?                      @      �?              �?                                                              �?      @     �Q@fffff�t@                                      6@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @     @3@������y@                      �?              O@      �?       @      �?       @       @       @       @       @       @       @              @�����|\@fffff�@                      �?      �?     �P@              �?               @       @       @       @       @               @              �?�����K@ffff�O�@      �?      �?                      �?      �?              �?                               @                                       @����̬R@����̬R@              �?                      0@      �?       @      �?                                       @       @              �?       @�����X@����̴�@      �?                              G@              �?                               @       @                      �?              �?������@@fffff�@      �?              �?              R@      �?       @                       @       @       @       @       @       @      �?      �?�����\U@    �S�@                                      J@      �?                                       @                       @              �?       @������M@fffffǧ@      �?              �?      �?      =@      �?       @                       @       @               @       @                      �?fffffT@�����G�@      �?                              *@      �?       @      �?       @                               @       @                      @������X@     9�@      �?              �?              7@      �?       @      �?               @       @                                               @     U@fffff��@      �?                      �?      6@      �?               @      �?      �?      �?      �?      �?      �?                      �?fffff&4@     {@                      �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@�����؇@      �?              �?              >@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?33333�4@�����X�@                      �?              R@      �?       @               @       @       @               @       @       @      �?      �?������T@����Y�@                      �?      �?      E@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @�����3@�����·@                                      5@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?������4@     4{@                      �?             �Q@      �?       @               @       @       @       @       @       @       @              �?33333SV@ffff���@      �?              �?      �?      9@      �?               @      �?      �?      �?      �?      �?      �?      �?               @������3@fffff�y@      �?      �?      �?             �B@      �?       @      �?                                       @       @              �?       @      W@�����"�@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@     `\@                      �?              A@      �?       @               @       @               @                                       @33333SO@�����š@                      �?              R@      �?       @      �?       @                                               @                �����T@�����i�@              �?                     �Q@      �?       @               @       @       @       @       @       @       @              @fffffvV@3333s��@                      �?      �?      @              �?                                                                              @�����9@     `_@      �?                              .@      �?       @                                                                               @fffff�I@     �@                      �?      �?     @Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ������9@�����%�@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�4@�����|c@              �?      �?             �M@      �?       @      �?       @       @       @       @                      �?      �?       @33333�W@ffff�k�@                      �?      �?      1@      �?       @                               @       @                      �?      �?      @������N@����̺�@                                     �B@      �?       @      �?       @       @       @                                                ������V@�����l�@                                     �L@              �?               @               @       @                      �?      �?      �?����̌D@    ���@      �?                              P@      �?       @      �?       @               @       @               @       @              �?     �X@3333s��@                      �?      �?      "@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y4@33333�g@      �?              �?      �?      (@      �?                                                       @                      �?      @fffff&L@33333��@              �?                     �J@      �?              �?               @                                              �?      �?33333sR@3333�G�@      �?              �?      �?     �E@      �?       @      �?                       @       @       @       @      �?      �?      �?33333Z@�����c�@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @              �?fffff\@3333��@      �?                              I@              �?               @                       @                      �?      �?      @33333�A@�����S�@                      �?              M@      �?                       @       @                       @                      �?      �?     PP@33333��@      �?      �?      �?             @P@      �?              �?                                                      �?      �?        ����̼Q@33333˱@                      �?              8@      �?       @      �?                       @                                      �?      @������S@�����"�@              �?      �?      �?     �Q@      �?       @               @       @                       @              �?               @�����LQ@    �v�@                      �?      �?     @P@      �?       @               @       @       @       @       @       @       @                33333�V@3333�K�@                                      $@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @������3@     �h@      �?              �?              E@      �?       @      �?                       @       @       @       @      �?      �?       @33333[@ffff&�@      �?                              >@      �?              �?               @                       @       @      �?      �?             @X@�������@                      �?              R@      �?       @               @               @       @       @       @       @      �?        �����9U@����L��@      �?              �?      �?     �E@      �?       @               @                       @               @      �?      �?      �?������Q@3333�ʨ@                                      R@      �?       @               @       @                                       @                     �M@     ��@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                       @33333�4@33333�4@              �?                      @      �?              �?                                       @       @              �?       @fffffVV@fffff��@                                      @              �?                                                                               @     @9@33333sM@                      �?              I@      �?       @      �?       @       @               @       @       @      �?               @33333#[@3333��@                                      2@      �?              �?               @       @                                               @33333sS@fffff:�@      �?              �?             �Q@      �?              �?       @       @       @       @               @       @              �?     @Y@    ���@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@33333#P@                                     �J@      �?       @      �?       @       @       @                                               @33333�V@333339�@      �?                             �L@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�4@fffff��@      �?                              8@      �?              �?               @       @       @                              �?       @�����|U@����Lv�@      �?                               @      �?                                                                                      @������F@     @T@                                       @      �?       @      �?                                                              �?      �?fffff�R@33333'�@      �?              �?              "@              �?                                       @       @                              @33333SD@33333�t@      �?              �?      �?      6@      �?                       @               @       @       @              �?      �?             �P@33333 �@      �?              �?      �?      R@      �?       @               @               @       @       @       @       @      �?      �?33333�T@����Lͷ@      �?                              9@      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff&4@�����@      �?      �?                      0@      �?       @      �?                                       @                      �?       @fffff�U@     �@                      �?      �?      .@      �?       @      �?               @       @               @       @              �?        fffffVZ@     ]�@                                      =@              �?                                                                      �?      �?�����9@�����F�@      �?      �?                      @      �?              �?               @                               @              �?       @33333cU@     �y@                      �?             �B@      �?       @                       @               @               @      �?              @fffffR@�����Ĥ@      �?                              @      �?       @                                                                               @33333�G@������k@                      �?      �?      5@      �?                               @                       @              �?      �?      �?�����lM@�������@      �?      �?                      &@      �?              �?                                               @              �?      �?������S@�����݉@      �?                              8@      �?       @               @                                                      �?        33333�K@33333�@      �?                              �?      �?                                                                                      @�����LF@�����LF@                      �?      �?     �N@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �3@fffff~�@                      �?              D@      �?       @                       @                       @              �?                33333�O@     ��@      �?              �?      �?     �K@      �?                       @                                       @      �?              �?������M@     ��@                                      3@      �?              �?       @               @       @       @       @              �?       @fffff�Z@�����9�@      �?              �?             �@@      �?       @      �?               @       @                       @              �?       @fffffVW@     (�@                                     �B@      �?       @               @                               @              �?                �����)P@3333�W�@                      �?      �?      9@      �?       @      �?                       @                       @              �?       @fffffFV@����̀�@                      �?              R@      �?       @      �?       @       @                                       @      �?        33333U@    @��@      �?              �?              F@      �?                       @       @               @                      �?      �?        ������M@ffff�W�@      �?                              Q@      �?       @      �?       @       @       @                       @       @      �?        fffff�Y@����Y�@      �?              �?              2@      �?       @      �?       @                               @       @              �?       @������X@�����;�@                                      @      �?                       @       @                                                       @����̬K@fffff�d@                      �?              $@      �?               @      �?      �?      �?      �?      �?      �?              �?        33333�3@     xg@      �?              �?             �Q@      �?       @               @               @       @               @       @      �?      �?33333�R@�����ô@      �?                               @      �?              �?                                               @              �?       @�����T@33333�f@      �?              �?             �H@      �?       @               @               @       @       @       @      �?               @fffffU@3333���@      �?                              2@      �?       @      �?               @                                              �?       @�����)T@�������@      �?              �?             @Q@      �?       @      �?       @       @       @       @       @       @       @      �?        33333#\@    �~�@                      �?              2@      �?              �?                       @               @       @              �?      �?������W@     F�@      �?                              @      �?       @                                       @       @                      �?      @     PP@�����<j@                                     �C@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�4@�����Ӈ@              �?      �?      �?      <@              �?                                               @                      �?       @33333�A@33333m�@      �?                              @      �?                                               @       @       @              �?       @fffffVQ@33333�g@                      �?      �?     �I@      �?              �?       @       @                                              �?        ������S@����e�@                      �?             �H@      �?       @                                                                      �?      �?33333J@    �/�@      �?                              �?      �?              �?                                                              �?       @fffffFQ@fffffFQ@      �?                              ,@      �?               @      �?      �?      �?      �?      �?      �?              �?       @�����4@����̴r@      �?      �?      �?               @      �?              �?                       @               @       @              �?      �?     �W@����̴f@                      �?               @      �?       @      �?                                               @              �?      �?�����LU@33333��@      �?                             �C@      �?                                               @                       @      �?        fffff�H@�����̞@                                      4@      �?                                                                              �?       @�����,F@33333��@                                     �F@      �?       @      �?                       @                       @              �?      �?33333SV@ffff&`�@      �?      �?      �?              @@      �?       @      �?               @       @               @       @                        fffff�Z@    ���@      �?              �?             �N@      �?       @      �?               @               @       @               @      �?       @fffff�W@����L�@                      �?             �I@              �?                       @                       @       @              �?       @33333�H@3333��@                      �?      �?     �J@              �?               @       @       @                       @              �?        �����YH@fffff~�@      �?              �?      �?      C@      �?       @               @               @       @       @       @       @      �?        �����YU@     ©@      �?                              "@      �?                       @               @       @       @                      �?      @     `Q@     j�@                      �?      �?      ,@      �?       @       @      �?      �?      �?      �?      �?      �?                      @����̌9@33333Gw@              �?                     �H@      �?       @      �?       @       @       @       @               @      �?                     �Y@33333.�@                                      �?      �?                       @                                                      �?        �����9H@�����9H@      �?                              �?      �?              �?                                                              �?      @33333�Q@33333�Q@      �?                             �F@      �?              �?       @       @       @       @       @       @      �?              �?�����\@����٧�@                                      @      �?       @      �?                                       @       @              �?      @�����yW@�����m~@              �?      �?             �G@      �?       @      �?       @                                                               @fffffT@3333��@      �?                              B@      �?                               @               @               @      �?      �?      @�����YP@����̄�@              �?      �?              L@      �?       @      �?                               @                              �?        fffff6S@    ���@                      �?      �?      6@      �?                               @                       @       @      �?      �?             `Q@�����h�@      �?              �?              ,@      �?       @      �?                                               @              �?       @�����IU@�����̑@                      �?      �?      3@      �?               @      �?      �?      �?      �?      �?      �?                      @3333334@33333�w@                      �?      �?      K@      �?       @               @       @       @       @       @       @       @              �?33333�V@     e�@                                      "@      �?              �?                                       @                      �?        �����iS@33333Q�@      �?      �?      �?      �?      J@      �?       @                       @       @               @       @      �?      �?       @fffff6T@����߯@      �?      �?      �?             �O@              �?               @                       @                      �?                �����B@�������@      �?      �?                      A@      �?              �?                                                                      �?�����IQ@33333ơ@                      �?      �?      L@      �?       @               @               @                       @      �?      �?             0Q@     ��@                                      @      �?       @      �?                                                                        ������R@������j@              �?      �?      �?      R@      �?       @               @       @       @       @       @       @       @      �?        ������V@3333s<�@      �?      �?      �?              >@      �?       @      �?                                                                      @�����yS@ffff�^�@                                      "@      �?              �?       @                                                      �?      �?     �R@33333��@                      �?      �?      ;@      �?       @       @      �?      �?      �?      �?      �?      �?       @               @     �8@�����χ@      �?              �?      �?      Q@      �?       @                       @               @               @       @              �?33333�Q@3333���@                      �?             �I@      �?              �?                                                                      @�����IQ@33333��@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�2@333333g@      �?                             �O@      �?              �?       @       @       @       @       @       @       @              �?�����L[@    ���@      �?                              �?      �?       @      �?               @                                              �?       @������S@������S@                      �?      �?      7@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?������9@     �@                      �?              Q@      �?       @      �?       @       @       @               @       @       @      �?        33333�[@�������@                      �?             �H@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?      3@�������@      �?              �?      �?      4@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@      y@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     �7@     =�@                      �?              .@      �?              �?       @               @               @       @                       @     pY@������@                      �?              R@      �?       @               @               @       @       @       @       @      �?      �?�����U@3333sз@              �?                      <@      �?       @      �?                       @       @       @       @              �?       @33333�Y@����L��@                                      @      �?       @      �?                                                                       @fffffS@�����p@      �?                              *@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@     �p@      �?      �?      �?              1@      �?              �?                                               @                             `T@�����Ĕ@              �?                       @      �?              �?                                                              �?       @������Q@33333�a@                      �?              P@              �?               @               @       @               @       @               @������G@     ��@      �?                             �C@      �?       @                                       @                       @      �?      �?������J@fffff1�@                                      :@      �?              �?                                                              �?      �?33333CQ@�����^�@                                      .@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@������t@                              �?      1@      �?                                                       @       @              �?      @�����,P@fffff�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      �?������3@������3@      �?                              (@      �?                               @               @                              �?      @     �J@33333E�@                                     �E@              �?                               @               @       @              �?        fffff�H@fffff8�@                      �?      �?      K@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����Y4@fffff�@      �?                              R@      �?               @      �?      �?      �?      �?      �?      �?       @                �����L3@33333�@      �?                              $@      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@�����!h@      �?              �?      �?     �P@      �?                       @               @       @                       @      �?        333333N@fffff�@                      �?             �J@      �?              �?       @       @       @       @       @       @      �?               @     �[@    �˶@      �?      �?                       @              �?                               @                                      �?       @ffffff=@����̼k@                      �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @                ������3@fffff��@                      �?              :@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @      :@fffff`�@      �?                             �J@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �����8@�����W�@      �?      �?      �?              9@      �?       @      �?       @                                       @      �?      �?       @33333CV@ffff��@      �?              �?             �F@      �?       @      �?               @                                                        �����YT@3333��@      �?              �?              �?              �?                                                                      �?       @33333s7@33333s7@      �?                             �L@      �?       @      �?                                       @              �?      �?       @������U@    @K�@      �?                              C@      �?                                       @       @               @      �?      �?      @fffff&O@�����e�@      �?                              ,@              �?                       @                                              �?      @�����?@33333;z@                                     �G@              �?               @               @       @                       @              @33333�D@     M�@              �?                      @      �?                                                                                       @     �F@fffff�_@                      �?      �?      1@      �?              �?                       @       @       @       @      �?                fffff�X@����̣�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@�����4@              �?      �?              >@      �?       @      �?               @                       @                      �?       @33333�V@fffff��@                      �?              .@      �?              �?               @                                                        fffff�R@33333j�@      �?              �?             �N@      �?       @      �?                                       @       @      �?      �?              X@3333�)�@      �?              �?              @      �?              �?                       @       @                              �?      @fffff&T@fffff�s@                                      2@      �?               @      �?      �?      �?      �?      �?      �?              �?      @����̌3@     Tx@      �?              �?      �?     �P@      �?       @      �?               @       @                              �?               @������U@������@              �?      �?              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @������4@������4@      �?                              2@      �?                       @                                                               @33333�H@fffffV�@      �?              �?      �?      �?      �?                                                                                       @fffffFF@fffffFF@      �?              �?              N@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@�������@      �?                               @      �?              �?               @                       @       @                       @������W@������d@                                      6@      �?       @               @                       @                              �?      @fffff�M@     ��@              �?      �?              4@      �?                               @                               @              �?       @      N@fffff��@                                      ?@              �?               @       @               @               @       @      �?        ������H@fffff��@      �?              �?              6@      �?               @      �?      �?      �?      �?      �?      �?              �?        33333s4@�����x}@      �?              �?      �?     �J@      �?       @                               @       @       @       @      �?      �?      @     �S@ffff�̮@      �?              �?      �?     �C@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @������7@fffff>�@      �?      �?                     �L@      �?                                       @       @                      �?      �?       @     �J@�������@              �?                      J@      �?       @      �?       @       @       @               @       @                      �?fffff[@����L϶@      �?              �?      �?      @@      �?              �?       @       @                               @      �?      �?       @33333�V@3333���@                      �?      �?     �Q@      �?       @      �?       @       @       @       @                       @                �����yW@������@      �?                             @Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333�7@fffffĚ@      �?              �?              2@      �?       @      �?                                       @       @              �?       @     �W@�����o�@      �?              �?      �?      R@      �?       @      �?               @       @       @       @       @       @      �?             \@ffff�i�@      �?      �?      �?              =@      �?       @      �?               @       @                       @              �?       @������W@fffffr�@                      �?              Q@      �?       @               @       @       @       @                       @              �?������Q@����Y/�@                                       @              �?                                                                               @     �8@333333G@      �?                              A@      �?       @      �?               @               @       @       @              �?       @fffffVZ@����L��@      �?                              I@      �?              �?       @       @               @               @              �?      �?     `W@    ���@                                       @      �?              �?                                               @                       @33333#T@33333g@                      �?              @      �?                                               @                              �?       @33333�H@������p@      �?                              @      �?              �?                       @       @       @                      �?      @fffffvV@fffff�n@                      �?             �Q@      �?                       @       @       @       @       @       @      �?      �?        333333U@������@                      �?      �?      R@      �?       @      �?               @       @       @               @       @      �?        ������X@3333sٻ@      �?                             �B@              �?               @       @               @                       @      �?      @fffffFD@fffff��@                                      2@      �?              �?                                                              �?       @fffff�Q@     �@      �?      �?                      8@      �?       @                       @                                                      �?ffffffK@33333-�@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                       @     @3@     @3@      �?                              @      �?                               @                                              �?       @����̬I@�����dp@                                      ,@      �?                       @                                                                �����I@     ,�@      �?      �?      �?             �H@      �?       @      �?       @       @       @                                      �?       @�����V@3333s?�@                              �?      �?      �?                       @                                                              @33333�H@33333�H@                      �?              =@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @����̌3@fffffN�@      �?                             �D@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff&4@������@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �3@fffff6X@      �?      �?      �?             �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @                      9@     w�@      �?                              D@              �?                       @               @                      �?              �?      B@�������@      �?              �?      �?      Q@              �?               @       @       @       @               @       @      �?      @333333L@ffff�خ@                      �?             �Q@              �?                       @       @       @       @       @       @                      M@ffff�1�@                      �?              A@      �?       @      �?                       @               @       @              �?       @�����Y@����L��@                                      C@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@     ,�@      �?                              (@              �?                       @               @                                      @      A@33333�{@                                      D@      �?       @      �?                                               @                        fffff�T@    ���@                      �?             �E@      �?                       @               @       @       @       @       @      �?       @33333�S@������@      �?              �?      �?     �C@      �?                       @       @       @                              �?               @fffff�M@3333�O�@                      �?              Q@      �?                       @                       @                      �?                33333�K@������@              �?                     �Q@      �?       @      �?       @       @               @       @              �?      �?      �?������X@    @�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff3@�����LI@      �?              �?              R@      �?       @      �?       @       @               @               @       @      �?        33333#Y@������@                              �?     �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?      9@fffffi�@      �?              �?      �?      O@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ������8@     �@      �?              �?      �?      @      �?                                                                              �?        �����LF@�����Lp@      �?      �?      �?              =@      �?       @      �?                               @                              �?       @33333�S@����ݢ@                      �?      �?       @              �?                                       @                                        �����=@     `F@      �?                      �?     �Q@      �?       @      �?       @               @               @       @       @                ����̬Z@    @ּ@                                     �D@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�4@33333�@                                       @      �?                               @                                                      @������H@������Y@      �?              �?      �?     �I@      �?       @      �?       @       @               @       @       @      �?              �?33333�[@fffff6�@                                       @      �?                               @               @                              �?      �?fffff�K@     �Y@                      �?              R@      �?       @               @       @       @       @       @       @       @                33333V@�����x�@                      �?      �?      @@      �?       @      �?       @                               @                               @ffffffV@�������@      �?                             �P@      �?              �?       @               @       @       @       @       @      �?        �����iZ@    ���@      �?      �?      �?             �Q@      �?              �?       @       @       @               @       @       @              �?fffffVZ@ffff�W�@      �?              �?             �M@      �?       @      �?                                               @      �?               @33333cU@ffff�ܳ@                      �?      �?     �D@      �?                       @                       @       @       @      �?      �?      �?����̬R@����L�@              �?                      @      �?              �?                       @                                              @33333�R@�����\i@      �?                      �?      C@      �?       @      �?                       @               @       @              �?             �X@����L��@      �?                               @      �?              �?                                                              �?      �?33333�Q@     �c@                                     �D@              �?                       @                               @              �?       @�����,D@fffff7�@      �?                              ?@      �?       @      �?               @                                              �?       @�����IT@������@                                      7@      �?       @      �?       @                               @                      �?        33333�V@������@      �?                              *@      �?                               @               @       @       @                      @fffffVR@fffff�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff&3@�����_@                                     �Q@              �?               @       @       @       @                       @      �?        �����LF@����L�@                                      $@      �?                                               @               @              �?      @�����yN@fffff��@                      �?      �?      P@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @fffff�8@     �@                                      �?      �?                               @                                                       @     �H@     �H@                                      �?      �?              �?                                               @              �?       @������S@������S@                      �?              (@              �?                               @               @       @              �?        ������H@33333I�@      �?      �?      �?              B@      �?       @      �?               @                       @       @              �?       @      X@33333ت@      �?              �?      �?      R@      �?              �?       @               @       @       @       @       @      �?      �?�����9Z@���̌��@      �?      �?                      $@      �?              �?                                               @              �?       @     �S@fffff̈@      �?      �?                      3@      �?       @      �?                       @                                      �?       @fffff�S@     ��@                      �?      �?      A@              �?               @               @       @       @       @      �?              @     �N@�����$�@                      �?      �?     �F@              �?                       @       @       @               @      �?                     �I@     ��@      �?              �?             �N@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?����̌4@     ��@                                     �M@      �?       @      �?       @       @       @                       @              �?        ������X@3333���@      �?      �?      �?              A@      �?       @      �?                                                              �?       @33333�R@������@              �?      �?              Q@      �?                               @       @       @                      �?      �?        33333SN@������@      �?                              @      �?              �?                       @                                      �?        33333�R@ffffft@      �?                      �?      @      �?              �?                                                                       @�����iQ@33333�k@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?        �����i\@    ���@      �?                              ;@      �?                       @               @       @       @       @      �?               @�����lT@����I�@      �?                               @      �?                               @               @       @                      �?       @������P@�����G�@                                      $@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�����L3@fffff&g@                      �?             @P@      �?       @      �?               @       @       @       @       @      �?      �?      �?33333[@ffff�λ@              �?      �?              @      �?              �?                                                                       @33333�Q@������r@      �?                              <@      �?              �?                       @       @               @                       @     �V@����L��@              �?      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?����̌3@33333ؖ@      �?                      �?      7@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@33333}@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @               @������\@�����N�@      �?              �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������4@������@                      �?      �?     �Q@      �?       @               @                                       @      �?                �����LP@ffff&��@                                      5@      �?                       @               @       @                      �?      �?       @      N@fffff��@      �?                              :@      �?       @               @       @                                      �?               @fffff�N@����̷�@      �?              �?      �?     @P@      �?       @      �?       @               @       @       @       @       @                �����)[@3333��@              �?      �?              K@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�2@fffff�@      �?              �?              R@      �?       @      �?       @       @       @               @       @       @      �?       @�����i[@    @Ⱦ@      �?              �?      �?       @      �?       @               @       @               @               @       @      �?      �?�����	S@fffff.�@                      �?      �?      &@              �?               @                                                      �?       @������=@33333�u@                      �?             �I@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �9@     �@                      �?      �?      Q@      �?       @      �?               @               @                      �?      �?        ������T@fffffe�@      �?                      �?      Q@      �?       @               @       @               @       @       @       @      �?             �U@    ���@      �?                      �?      &@      �?       @      �?                       @                                      �?      @     �S@fffff��@      �?                               @              �?                               @               @       @              �?       @     �H@fffff�V@                                      @      �?              �?                                                              �?        ������Q@     q@                      �?      �?      P@      �?       @                       @                                      �?      �?        ������J@3333���@                                     �K@      �?       @      �?                                                              �?       @fffffFR@ffff�0�@                                     �I@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�4@     �@      �?              �?      �?      (@      �?               @      �?      �?      �?      �?      �?      �?              �?       @fffff&5@����� s@      �?              �?              R@      �?       @      �?       @               @       @       @       @       @      �?      �?������[@������@                                      M@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����Y8@fffff?�@              �?                      D@              �?               @       @                       @       @              �?       @fffff�K@3333�z�@      �?              �?      �?     �O@      �?       @      �?               @       @               @       @       @      �?        333333Z@    @Ź@      �?      �?      �?              8@      �?              �?                       @               @       @              �?       @�����IW@����n�@                      �?             �N@      �?       @      �?                       @       @       @       @      �?      �?        33333�Y@����Yv�@      �?              �?              @      �?       @      �?                                                              �?       @������R@fffff�r@      �?              �?              R@      �?              �?                       @               @       @              �?       @������W@����Y[�@                              �?      �?      �?                       @       @               @                              �?       @      N@      N@      �?                      �?      "@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@     �g@      �?              �?      �?      K@      �?       @                       @               @       @              �?      �?       @����̬Q@     t�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����3@�����3@      �?              �?      �?      A@              �?                                       @       @               @      �?       @fffffFD@fffff��@      �?                              @      �?                                                       @                      �?       @333333L@33333[m@      �?      �?                     �G@      �?       @                       @               @                       @                ������M@     ��@              �?                       @      �?       @      �?               @       @               @       @              �?       @     `Z@fffff�@                                      <@      �?                       @       @                                                       @fffffL@�����ʗ@              �?                      ,@              �?                                               @       @              �?       @�����,G@������@      �?              �?             �P@      �?       @      �?       @               @               @       @       @      �?      �?33333�Z@����YE�@      �?                              @      �?                                                       @                              @�����lK@fffff&w@                                      6@      �?              �?       @                       @               @              �?       @33333CV@     y�@                                      "@      �?               @      �?      �?      �?      �?      �?      �?                        fffff&4@������m@                      �?      �?      "@      �?                       @       @       @       @                                      @     @P@fffff��@      �?              �?      �?     �D@      �?       @                       @       @               @              �?                      Q@ffff�/�@      �?              �?      �?     �B@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@fffff(�@      �?                              $@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?      4@33333�h@                      �?             �Q@      �?       @      �?                       @               @       @      �?      �?       @     pY@����L��@      �?              �?              O@      �?                               @       @       @                       @      �?      �?33333N@fffffR�@      �?                              @      �?              �?                                                              �?      @ffffffQ@������i@                      �?              9@              �?                                               @                      �?              A@     ��@              �?      �?              9@      �?              �?               @       @                       @                        �����V@����L�@      �?              �?              R@      �?       @               @       @       @       @                       @              @�����	Q@3333�Ȳ@                      �?      �?      R@      �?       @      �?       @                                               @                33333�S@3333�b�@                              �?      2@      �?       @               @                                                              @33333�L@������@              �?                     �P@      �?       @                       @                                                       @33333sK@     �@      �?              �?             �L@              �?                       @       @       @       @       @       @      �?             �L@ffff惩@              �?                      1@      �?       @      �?                                       @       @              �?       @����̌W@����� �@                      �?             �O@      �?       @      �?               @                                              �?        33333cT@������@                                      2@      �?              �?                                                              �?       @33333sQ@������@              �?      �?             �Q@      �?       @      �?       @       @       @       @       @       @       @      �?       @�����i\@ffff�"�@      �?                              L@      �?                               @       @       @       @       @       @      �?      �?33333sT@3333s��@                                      (@      �?              �?               @                               @              �?       @fffff&U@�����ʏ@      �?              �?      �?       @      �?              �?       @                               @       @                       @fffffFX@�����g@                                      7@      �?               @      �?      �?      �?      �?      �?      �?              �?      @     �3@33333c}@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333s3@33333s3@      �?      �?                     �P@      �?       @      �?                                                              �?      @������R@�����ĳ@                      �?      �?      @      �?              �?                                       @                      �?      @������S@     �r@      �?              �?      �?      Q@      �?       @      �?               @                       @       @      �?      �?      �?33333CY@    �r�@      �?              �?      �?     �Q@      �?              �?       @       @       @       @       @               @      �?      �?fffffFY@�����R�@      �?      �?      �?             �K@      �?       @               @       @                                      �?              �?      N@33333�@                                      .@      �?       @      �?               @                                              �?       @     �S@fffff_�@              �?                      $@              �?                                                       @              �?       @�����YA@����̜t@      �?                              @              �?                                       @                                       @ffffff>@������T@              �?      �?             �Q@      �?       @      �?                                                       @      �?      �?������R@fffff#�@      �?      �?                      ,@      �?              �?                                       @       @                      �?����̜V@fffffȓ@      �?      �?      �?              "@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@������f@      �?              �?      �?      $@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333s4@�����Ln@                      �?      �?     @Q@      �?       @      �?       @               @                              �?                �����U@�����ض@      �?              �?      �?     �L@      �?                       @       @               @                      �?              @������M@�����j�@                      �?              2@              �?                               @               @                      �?       @fffff�C@������@                      �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@�����s�@      �?                      �?      �?              �?                       @                                              �?      @�����Y?@�����Y?@                      �?      �?      8@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�����5@fffff�~@      �?                              �?      �?              �?                                                              �?       @fffffVQ@fffffVQ@      �?                      �?       @      �?               @      �?      �?      �?      �?      �?      �?                        33333s3@fffff�c@                      �?      �?      M@      �?                                                                      �?      �?      @�����F@����ڢ@      �?              �?              @      �?              �?                       @               @       @              �?       @����̜W@�����!@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@     `S@      �?              �?             �Q@      �?       @               @       @       @       @       @       @       @                33333�V@     �@      �?                      �?      @      �?                                                       @                      �?      �?�����YK@fffff.e@      �?              �?      �?      O@      �?       @      �?                       @               @               @      �?      �?fffffFV@ffff�#�@      �?              �?      �?     �P@      �?                       @       @       @               @       @       @              �?fffffVT@������@      �?                              D@      �?       @      �?                       @       @       @       @                        333333Z@3333�#�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @������4@������4@      �?      �?                      P@      �?       @      �?       @       @                       @       @              �?             �Y@ffff���@                      �?              R@              �?               @       @       @                       @       @      �?       @������H@ffff���@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?             @3@     @3@      �?              �?             �O@      �?              �?       @       @       @       @       @       @       @      �?      �?fffff�[@3333�1�@                                      �?      �?              �?                                                              �?       @     �Q@     �Q@      �?                              @      �?       @      �?               @       @                                      �?       @33333SU@fffff�z@                                      Q@      �?                       @               @                              �?      �?      �?�����9K@ffff浬@      �?      �?      �?      �?     �P@      �?       @      �?                       @               @       @              �?      �?     �X@ffff&��@      �?                             �O@      �?       @      �?               @       @               @       @       @      �?             0Z@    ���@      �?              �?             �Q@      �?              �?               @       @       @       @       @       @      �?       @     PZ@    �{�@      �?              �?              8@      �?       @               @                       @                      �?      �?       @�����,M@������@      �?                              Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        fffff&8@fffffk�@              �?      �?      �?     �Q@      �?       @      �?               @       @       @       @       @      �?      �?       @������Z@�����3�@      �?              �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?             �\@ffff��@                      �?              R@      �?       @      �?       @       @       @       @       @               @      �?        ������Y@ffff愽@              �?                      @      �?       @                                                                              @     `H@33333{f@      �?      �?                      K@              �?                       @       @               @       @      �?      �?       @������K@ffff�-�@      �?                      �?      P@      �?              �?               @               @       @       @              �?      �?������X@33333�@              �?      �?              @      �?       @      �?               @                                              �?       @     @T@fffff:w@      �?              �?      �?     �P@      �?       @      �?               @       @               @       @      �?      �?       @�����YZ@3333sM�@              �?                      &@      �?              �?                                       @       @                        �����lV@�����^�@      �?              �?      �?     �P@      �?       @      �?               @                               @              �?        33333cV@�����@      �?                              7@      �?                                                       @       @      �?      �?        �����9P@33333��@                      �?              P@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333s3@fffff�@      �?              �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?����̌4@fffff�@                                      4@      �?       @      �?       @                               @                      �?        fffffFV@     ]�@      �?                              *@      �?              �?                                                              �?       @������Q@     �@                              �?      0@      �?              �?                                       @                      �?       @     @T@�������@      �?                               @      �?                       @               @                                      �?      @����̌K@fffffV\@      �?                             �A@      �?               @      �?      �?      �?      �?      �?      �?       @              @     @3@33333/�@      �?                              &@      �?              �?                       @                       @                       @333333U@     Ƌ@      �?                      �?      *@      �?                                                                                      @      F@����̚�@      �?      �?      �?               @      �?                                       @       @               @              �?      �?�����P@�����-�@      �?                              <@      �?              �?               @               @       @              �?      �?             �V@����Lg�@                                      I@      �?              �?               @               @       @       @       @      �?      @�����Y@3333s��@                      �?              ?@      �?              �?               @                               @              �?        fffff�T@����L�@      �?              �?              @      �?              �?                                                              �?       @fffffVQ@�����1|@                      �?      �?      C@      �?                       @       @                                                       @     @K@����8�@              �?      �?              @@      �?       @      �?                       @                                              @33333�S@     �@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              �?����̌3@333333Q@      �?              �?             �D@      �?       @                               @               @       @      �?      �?       @     @R@fffffr�@      �?              �?             @P@      �?       @               @               @       @               @       @                �����	S@���̌A�@      �?              �?              C@              �?               @       @               @       @       @       @      �?              N@fffff"�@      �?              �?      �?     �Q@      �?       @      �?               @               @                       @      �?       @333333U@fffff�@                                       @      �?              �?                                       @       @              �?       @������V@fffffe@      �?              �?      �?     �K@      �?       @      �?                       @               @                      �?      �?������V@ffff&�@      �?              �?      �?      @      �?              �?       @       @                       @                               @fffffvV@�����o@                      �?      �?      D@              �?                       @                       @       @              �?       @�����lI@33333ҟ@                      �?      �?      >@      �?                                       @       @       @              �?      �?       @      P@������@      �?      �?                      �?      �?              �?                                                              �?       @�����iQ@�����iQ@      �?              �?              R@      �?       @      �?               @       @       @       @       @       @      �?      �?     p[@ffff�N�@      �?      �?                      @      �?       @      �?               @                                              �?       @fffffVT@fffff6m@      �?                              �?      �?              �?                       @               @                      �?       @fffff6U@fffff6U@                                      K@      �?              �?       @       @                       @       @      �?      �?      �?33333Y@ffff���@      �?                              @      �?                       @               @       @       @       @                      �?������S@�����4~@                                      �?              �?               @                                                              @fffff�=@fffff�=@      �?      �?      �?              (@      �?              �?                                               @              �?       @�����T@�������@                                      �?      �?                       @                                                      �?      �?�����LH@�����LH@                                     �J@      �?              �?               @       @               @       @      �?      �?      @33333Y@�����P�@      �?                             �D@      �?       @      �?               @       @               @       @              �?       @�����,Z@fffff��@      �?      �?      �?              R@      �?       @      �?       @       @       @               @       @       @      �?        33333c[@3333��@      �?                              @              �?               @       @       @       @                              �?      @     �E@     `k@      �?              �?              K@      �?       @      �?               @       @               @       @              �?       @33333Z@ffff&��@                      �?      �?     �P@      �?       @                               @       @               @       @      �?        �����yQ@ffff��@      �?                             �I@      �?       @               @                       @                      �?              �?33333�M@33333ǧ@      �?                              R@      �?       @      �?               @       @               @       @       @      �?       @������Y@�����ҽ@      �?                             �H@      �?       @      �?               @       @               @       @              �?        ������Y@����L��@      �?      �?                      2@      �?       @      �?                                       @       @              �?       @������W@33333b�@      �?      �?      �?             �@@              �?                       @       @       @       @                      �?       @      I@fffff[�@      �?                      �?      .@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @������8@fffffBt@      �?      �?      �?              @@      �?       @      �?               @       @                       @              �?       @     `W@�����5�@                                      G@      �?               @      �?      �?      �?      �?      �?      �?       @      �?       @�����5@�����H�@      �?              �?      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?      �?              @ffffff3@fffff��@              �?                      �?              �?                                               @                      �?       @�����9B@�����9B@                      �?      �?      Q@      �?       @      �?               @       @                               @      �?      �?�����U@    �r�@                      �?      �?      H@      �?                       @               @       @       @              �?                �����lQ@����L��@                      �?      �?      0@      �?                       @       @               @               @       @                     Q@fffffk�@                                      "@      �?              �?                                       @       @              �?        33333�V@     N�@      �?                              .@      �?              �?                       @               @                               @33333SU@fffff�@                      �?              O@      �?       @               @       @               @       @       @       @      �?       @�����<U@���̌�@      �?              �?              P@      �?              �?               @       @       @       @       @      �?      �?      �?����̜Y@������@                      �?      �?      O@      �?       @      �?               @               @       @       @      �?      �?      �?33333�Z@    �/�@      �?                              :@              �?               @                       @       @       @      �?              �?fffffFK@fffffK�@                                      K@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@�����ݐ@      �?                              @      �?       @      �?                                                              �?       @������R@������l@      �?                      �?      .@      �?                                       @       @                      �?              �?������K@fffff�@      �?                             �I@              �?               @                       @               @              �?      �?�����9F@�����@      �?                              ;@      �?                       @               @       @       @              �?              �?fffffVQ@33333�@      �?                              �?      �?              �?                                               @              �?       @     �S@     �S@      �?              �?      �?      C@      �?       @      �?               @       @               @                      �?       @������W@�����P�@                                      9@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?3333333@����̠�@                                      O@      �?                       @                       @               @       @      �?      @fffffFP@    ��@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?      �?              �?fffff�3@fffff>c@                      �?      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����4@�������@      �?              �?      �?     �P@      �?              �?       @       @       @               @       @      �?      �?        ������Y@����Lw�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����L3@�����L<@      �?                      �?      (@      �?               @      �?      �?      �?      �?      �?      �?       @                �����Y3@������j@      �?              �?             �E@      �?              �?       @       @       @                                      �?      �?fffff�U@����L��@                                      @      �?       @                                       @       @                      �?      @�����P@     �o@      �?      �?      �?              N@      �?              �?               @       @               @       @      �?      �?       @�����|X@     �@              �?      �?             @P@      �?       @      �?       @       @       @               @       @              �?      �?�����Y[@3333s;�@                      �?      �?      4@      �?       @      �?               @       @               @       @              �?        fffffvZ@����L�@                      �?      �?      P@      �?       @      �?               @       @                       @      �?      �?       @fffff6W@    �\�@                      �?      �?      P@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������3@������@      �?              �?              A@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����4@     8�@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?       @      5@      5@                                      1@      �?               @      �?      �?      �?      �?      �?      �?      �?                fffff�3@fffff2t@      �?      �?      �?              R@              �?               @       @       @       @       @       @       @      �?      �?�����<P@     ±@                                      @      �?       @      �?       @                                                      �?       @33333�S@     ({@                      �?             �J@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������4@fffff�@      �?                              =@              �?                                                              �?      �?      @������8@fffff��@      �?                              �?      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @      9@      9@                              �?     @P@              �?                       @               @       @               @              @     �F@ffff��@      �?      �?      �?              >@      �?       @      �?                               @       @       @              �?       @     `Y@����L˦@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @      :@     ��@      �?              �?             �D@      �?               @      �?      �?      �?      �?      �?      �?       @      �?       @     �3@������@                              �?     �A@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�����4@     $�@      �?                              F@      �?              �?                                                                      �?fffff6Q@ffff��@                      �?              8@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?ffffff4@�����,~@      �?                              J@      �?       @      �?       @               @       @       @       @       @      �?       @33333S[@fffffc�@      �?                              ;@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����Y4@����̜�@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @       @                ������\@�����N�@      �?              �?             �N@      �?                       @       @               @       @       @       @      �?      @33333CT@ffff���@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�4@fffff�4@      �?      �?      �?             @Q@      �?       @      �?               @       @       @       @       @       @      �?       @�����|[@    @ҽ@                                     �@@      �?       @      �?       @                                       @              �?       @������V@33333[�@      �?              �?      �?      "@              �?                       @                                              �?       @33333�=@fffffo@                      �?              5@      �?                       @               @       @       @       @      �?              @�����9T@�����˚@                                       @      �?               @      �?      �?      �?      �?      �?      �?       @              @     @4@������e@                      �?             @Q@      �?              �?       @       @               @       @       @      �?      �?      �?������Z@ffff�S�@                      �?      �?      R@      �?                       @       @       @       @               @       @      �?       @fffff�R@fffffu�@                      �?      �?     �D@      �?       @               @       @       @               @              �?      �?      �?fffff�S@fffff�@      �?              �?             �K@      �?       @      �?       @       @                       @                      �?       @     0X@ffff�v�@                      �?              H@              �?               @               @                       @              �?        fffff�F@      @              �?      �?              A@      �?       @      �?               @       @                       @              �?       @     �W@����#�@      �?      �?      �?              �?      �?       @      �?                                                                       @33333�R@33333�R@                                     �D@      �?              �?               @               @       @       @       @      �?        33333�X@����L�@                                      C@      �?       @                       @               @               @                      �?�����	Q@�������@                      �?      �?     @P@      �?       @      �?               @       @       @       @       @       @      �?      �?33333�[@ffff�M�@                      �?      �?      R@      �?       @               @       @       @       @       @       @       @                �����)W@     M�@                                     �N@      �?       @               @       @       @       @       @       @       @               @�����iV@3333���@      �?                              ?@      �?       @                       @               @       @                      �?       @33333�Q@����L�@                                      H@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ����̌8@�����ϒ@              �?                      2@      �?              �?               @                                              �?       @����̬R@fffff:�@                      �?      �?     �F@      �?                               @               @                      �?      �?      �?33333K@������@      �?                              "@      �?              �?                                                                      @33333�Q@     ��@              �?      �?              N@      �?       @      �?       @       @       @       @       @       @       @      �?        33333]@ffff��@      �?              �?      �?     @Q@      �?                       @       @               @       @       @       @                �����)T@���̌��@                                     �E@      �?       @      �?               @       @               @       @       @      �?       @fffff&Z@����ٗ�@      �?              �?      �?     �Q@      �?                       @       @       @       @       @       @       @                �����\U@ffff捷@                                      �?      �?              �?       @                                                              @33333�R@33333�R@                              �?     �E@      �?              �?       @       @               @       @       @      �?      �?      �?     �Z@����L��@      �?              �?              Q@              �?               @               @               @       @       @      �?        �����K@     ��@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @fffff�3@33333�d@      �?              �?      �?     �B@      �?       @               @               @       @                       @      �?      �?ffffffO@    �͡@      �?                              H@      �?       @      �?               @       @               @       @      �?      �?      �?fffff�Z@�����ڳ@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              @�����3@      J@                                      K@      �?       @      �?               @       @               @              �?      �?             �W@    ��@                      �?      �?      ?@      �?       @                       @               @       @       @       @                33333#T@33333O�@                      �?      �?      >@      �?       @      �?                       @               @       @              �?       @33333Y@����Ļ@                      �?      �?     @P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?      :@fffffۙ@                      �?               @      �?       @      �?                       @       @       @       @              �?       @�����Z@�����Yn@                      �?              Q@      �?       @               @       @       @       @       @       @       @      �?       @������V@3333��@                                     �@@      �?              �?               @               @                      �?      �?        ������S@3333���@      �?                             @P@      �?       @      �?       @                       @               @      �?               @33333cW@    @��@                      �?      �?     �P@      �?                       @                               @               @      �?       @     �M@�����9�@                      �?              &@      �?       @      �?       @                       @       @                      �?      �?�����X@33333�@                      �?      �?     �O@      �?                       @       @       @       @       @               @              �?33333�R@�����c�@      �?              �?      �?     �K@      �?              �?               @               @                                       @������S@3333s��@                                      A@      �?                       @       @                                      �?              @     �K@�����t�@                      �?      �?     �Q@      �?       @               @       @       @       @       @               @                ������S@����Lo�@      �?              �?              @              �?                                                                              @      9@     �S@      �?              �?             �O@      �?       @                       @               @               @       @              @     �P@ffff&��@              �?                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@������V@      �?                              @              �?                               @               @                      �?      @33333D@     X`@                      �?      �?      M@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����L4@     #�@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @      �?      �?������V@ffff�ֹ@      �?              �?      �?      B@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333s3@     ��@              �?      �?              R@      �?       @      �?       @               @       @       @       @       @      �?      @     p[@����Y��@      �?              �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     @8@������@                      �?      �?      R@              �?               @               @               @       @       @      �?      �?fffff�J@ffff��@                                      .@      �?       @                                                                      �?       @����̌H@fffff<�@              �?                      E@      �?       @      �?                                       @                      �?       @�����)U@3333���@      �?                      �?      �?      �?       @      �?                                       @       @              �?       @33333SW@33333SW@      �?              �?              R@      �?       @               @       @       @       @               @       @      �?        33333�T@���̌\�@      �?              �?      �?      "@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@����̬h@                      �?      �?     @Q@      �?       @               @       @               @       @              �?              �?�����lR@������@      �?              �?              E@              �?               @                               @                      �?        33333D@33333h�@              �?                      P@      �?                       @       @               @       @               @      �?      �?����̌Q@     ��@              �?                      R@      �?       @      �?               @       @       @       @       @       @               @������[@3333s�@                                      :@              �?                               @               @       @              �?      �?�����,I@     ��@      �?      �?                      �?      �?              �?                                       @                      �?       @fffff�S@fffff�S@      �?              �?      �?      G@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �3@     Ċ@      �?              �?      �?      @      �?       @      �?               @       @                                      �?        333333U@fffff>w@                                      O@      �?       @      �?       @       @       @                              �?      �?       @33333W@�����{�@      �?              �?      �?      @      �?                                                                                       @     `F@fffff�t@                      �?             �J@      �?              �?                       @               @       @      �?      �?        fffff�W@33333��@                      �?               @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@������D@      �?              �?              J@      �?       @               @       @       @       @               @      �?      �?      �?�����YT@3333s�@                              �?      �?      �?              �?                                               @                       @������S@������S@      �?                              *@      �?              �?       @                                                      �?      �?     pR@33333�@      �?              �?      �?      M@      �?       @      �?                                       @               @                     �T@����ܲ@                      �?      �?      R@      �?       @      �?       @               @       @       @       @       @              @������Z@3333���@      �?              �?             �E@      �?              �?       @               @       @                      �?      �?             U@    ���@      �?                              8@      �?       @      �?               @                       @       @              �?        ������X@3333�ɢ@      �?                              @      �?              �?                                       @                               @     �S@������p@                                      7@      �?       @               @                                                               @333333K@     ��@              �?      �?      �?      @      �?                                                                                       @      G@33333�f@      �?              �?      �?     �I@              �?               @       @       @               @       @      �?               @fffff�M@����L��@      �?                             �Q@      �?       @      �?                       @       @                       @      �?      �?������U@     �@      �?      �?      �?             @P@      �?       @      �?       @       @                       @               @      �?      �?�����,W@fffffP�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @     �3@     �3@                      �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?                      �?�����5@     xa@                                      �?      �?                                                       @                      �?       @33333SK@33333SK@                      �?              @      �?              �?       @               @                       @              �?      @�����9V@fffffb|@      �?                              *@      �?              �?               @       @                                      �?       @33333�S@�����k�@              �?                      ,@      �?       @      �?               @       @               @       @              �?       @fffff6Z@������@                                      0@      �?              �?               @                                                        fffff�R@fffff�@      �?              �?              G@      �?       @      �?               @       @               @              �?      �?       @������W@    �ذ@                                     �I@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ������3@�����'�@      �?                      �?      >@              �?                                               @       @              �?       @     @F@33333o�@      �?              �?              O@      �?       @      �?                       @       @       @       @       @      �?        fffff�Z@3333� �@      �?                              &@              �?                       @               @                              �?       @33333�A@������z@      �?              �?      �?      D@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     @9@33333w�@                                     �A@      �?              �?                       @       @       @       @      �?      �?       @     �X@     ��@                      �?              I@      �?       @      �?       @       @               @       @       @              �?        �����i[@������@                      �?      �?     �K@      �?       @               @               @       @       @       @       @      �?        fffffFU@3333�1�@              �?      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?     �\@�����}�@      �?                               @      �?       @                       @                                              �?      @333333K@fffff�\@      �?                              3@      �?                                       @       @                              �?      �?     �K@     Z�@                      �?      �?      �?      �?                                       @                                              @�����9I@�����9I@                                      @      �?              �?                                                              �?       @     �Q@fffff�l@                      �?      �?      @      �?              �?               @                               @              �?       @fffff�T@33333Cy@                      �?      �?     �G@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@33333��@                      �?      �?      L@      �?       @               @                               @              �?                �����LP@����Lp�@                      �?              K@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����4@�����9�@      �?                              K@      �?               @      �?      �?      �?      �?      �?      �?       @              @      4@�������@      �?              �?             �Q@      �?       @               @       @       @       @               @       @              �?�����T@ffff&_�@      �?                              3@      �?       @                                               @       @                      @ffffffQ@33333ʕ@                                      *@      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����L4@fffff6q@                                      7@      �?              �?       @                                                      �?             �R@     ʛ@                                       @      �?              �?       @       @                       @                      �?       @������V@     e@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@     �M@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     @3@     @3@      �?              �?              1@      �?              �?                       @               @       @      �?      �?        �����)X@     ј@      �?              �?              R@      �?       @               @       @       @       @       @       @       @      �?      �?�����,V@3333���@      �?              �?              @      �?                                       @       @                              �?      @fffff�K@�����Qc@      �?                              @      �?       @      �?               @       @               @       @                       @33333SZ@�����4�@      �?      �?                      O@      �?       @      �?               @       @       @       @       @      �?      �?             �[@����Y��@      �?                      �?      =@      �?       @      �?               @       @       @               @      �?              �?33333#Y@ffff��@                                      �?      �?                               @                                              �?       @�����LH@�����LH@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @������2@������2@      �?                               @      �?              �?                                                              �?      �?33333sQ@fffff�`@                                      *@      �?       @      �?                                               @              �?       @fffff&U@�����l�@                                      $@              �?                       @               @                                       @      B@     `w@      �?      �?                     �L@      �?       @                       @       @               @       @       @      �?             �S@33333V�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@�����Q@      �?              �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @              �?      4@�����x�@      �?              �?              ?@      �?       @                               @       @       @       @      �?      �?      @33333�S@     h�@      �?                              ?@      �?                                       @       @                              �?       @     �K@�����Κ@      �?              �?      �?      1@              �?               @               @               @              �?              �?�����9F@33333��@      �?              �?             �I@      �?       @      �?               @       @               @       @      �?      �?        33333�Z@�����z�@      �?                             �J@      �?              �?               @               @                              �?      @fffff&T@������@                      �?              4@      �?              �?                       @       @                              �?      @     @T@�����N�@                                      M@      �?                       @       @       @       @                       @      �?      �?�����9P@ffff榭@      �?              �?              9@      �?              �?                               @       @       @              �?      �?������W@3333�D�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @������3@������3@              �?      �?             �B@      �?              �?                       @       @       @                               @     �V@    �W�@      �?              �?      �?     @Q@      �?                       @       @       @                               @      �?             �M@�����˯@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@33333�T@      �?      �?      �?              �?      �?       @      �?                                       @                      �?       @33333�U@33333�U@      �?                      �?     �Q@      �?                       @       @       @       @       @               @      �?      �?�����9S@3333���@                                     �L@      �?       @      �?       @       @       @               @       @       @      �?        �����<\@     A�@                                      0@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����Y3@�����xr@      �?      �?      �?              F@      �?       @      �?                       @               @                      �?       @�����LV@fffff��@                                      9@      �?               @      �?      �?      �?      �?      �?      �?                      @�����3@������|@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@     �4@                                       @      �?              �?                                               @                       @     0T@fffff�c@      �?              �?      �?      1@      �?       @      �?                                       @       @              �?       @33333#W@fffff��@                      �?      �?      M@      �?       @               @               @       @       @               @              @33333�R@    �?�@                      �?             �N@      �?       @      �?               @               @               @       @      �?        fffff�W@     G�@                      �?             �B@      �?       @      �?                       @                                      �?      �?����̼S@����L/�@              �?                     �B@      �?       @      �?                                                              �?       @     S@����3�@                                      @      �?       @      �?                                                              �?       @fffff�R@33333��@                                     �A@      �?       @      �?               @               @                                      �?33333SU@     ˦@                      �?      �?     @Q@      �?       @      �?       @       @       @       @       @              �?      �?      �?fffffFZ@�����B�@                      �?              @      �?       @      �?               @       @               @       @              �?       @33333SZ@�����	�@      �?      �?                     �C@      �?       @      �?               @                               @                       @����̬V@    ���@                                      .@      �?              �?       @       @                       @       @              �?      �?fffff�X@�����I�@      �?      �?                      (@      �?       @      �?                       @               @       @              �?       @������X@�������@      �?                              .@      �?       @      �?       @                               @       @              �?       @������X@     {�@                      �?      �?     @P@      �?       @               @       @       @       @       @       @       @      �?      @����̜V@ffff�E�@                      �?      �?     �Q@      �?                       @               @       @       @       @       @      �?      �?     �T@�����o�@      �?                              @      �?       @      �?                       @               @       @              �?        33333cY@������r@      �?              �?      �?      Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �9@�����X�@      �?      �?                     �@@      �?       @      �?               @       @                                      �?      �?fffff�T@�����8�@      �?                              @      �?                                       @       @       @                                33333P@33333�{@      �?                             �A@      �?              �?               @       @               @       @      �?      �?        fffff�Y@33333T�@                      �?      �?      J@      �?       @      �?       @       @       @                       @                        ������X@fffff��@                      �?      �?      G@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�3@�������@      �?              �?             �F@      �?       @      �?               @       @               @       @              �?             �Z@������@      �?                              @              �?                                                              �?      �?      �?�����Y8@33333�b@                                      �?      �?              �?                       @                                               @33333�R@33333�R@                                      �?      �?              �?                                                              �?       @     `Q@     `Q@      �?              �?      �?      Q@      �?                       @       @       @       @                       @              �?33333SO@������@                      �?      �?      $@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����:@�����1l@      �?              �?      �?      N@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        33333�4@33333ړ@      �?              �?      �?      @      �?                                       @                                               @�����YH@     Du@                      �?      �?      K@      �?       @                       @       @                               @      �?        fffff�M@ffff�\�@      �?              �?             �Q@      �?                       @       @               @               @       @              @������P@ffff&8�@      �?              �?      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        33333s3@     @                      �?              =@      �?               @      �?      �?      �?      �?      �?      �?                      @������3@fffff�@                      �?      �?      B@      �?       @      �?               @       @               @                      �?        fffffVX@������@      �?              �?      �?      (@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @ffffff:@33333�s@      �?                             �K@      �?       @      �?                                       @       @              �?       @333333X@3333�@                                      &@      �?              �?       @                                                               @�����S@�����5�@              �?                      6@      �?              �?       @       @                                                       @�����lT@�����s�@      �?              �?      �?      J@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?������4@fffff��@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@����̬N@                      �?      �?      L@      �?       @      �?                       @               @       @      �?      �?      �?33333�X@3333s��@                                      O@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?������9@�����o�@                                      @      �?       @      �?                       @               @       @              �?       @      Y@     �@      �?      �?      �?             @P@      �?       @      �?               @       @               @       @      �?      �?        ������Y@3333s��@      �?                              ,@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?������8@33333t@      �?              �?              E@      �?       @      �?               @       @       @               @              �?       @������X@����*�@      �?              �?              9@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        33333�4@fffff�~@      �?      �?                      4@      �?       @      �?                                       @                      �?       @fffffU@�����D�@      �?      �?                       @      �?              �?                                                              �?       @�����lQ@������@      �?                      �?     @Q@      �?       @               @       @       @       @       @               @      �?      �?������S@���̌~�@      �?              �?              J@      �?              �?       @                               @                               @fffffU@ffff���@      �?              �?              P@      �?              �?       @                                                      �?      @33333cR@     ��@      �?                             �P@              �?               @                       @       @               @               @33333�E@fffff2�@      �?                              K@      �?                       @       @               @       @                      �?      @�����yQ@�����V�@      �?              �?      �?      &@      �?               @      �?      �?      �?      �?      �?      �?                        33333�4@������p@      �?              �?      �?      M@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @����̌3@33333S�@                                      "@      �?       @      �?                                               @              �?       @33333�T@fffff�@                                      @      �?       @      �?                                                                       @33333�R@fffff�y@      �?                              2@      �?       @      �?                                       @                                33333U@������@      �?              �?      �?      @      �?       @                                                                      �?       @33333sI@333333l@      �?              �?      �?      *@      �?       @                       @       @       @       @                      �?       @333333R@fffff�@              �?      �?             �E@              �?                       @       @               @       @                      �?fffff�K@fffffL�@      �?                              @      �?              �?                                               @                      @     �S@������z@                                      N@      �?              �?       @               @       @       @       @              �?        �����<Z@    �\�@      �?      �?      �?              >@      �?                               @                                              �?        333333I@     ޗ@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@     @_@                      �?             �Q@      �?       @      �?                       @               @       @      �?      �?       @�����iX@    �F�@      �?              �?      �?      I@      �?                                                                      �?      �?        ffffffF@3333�m�@      �?              �?              G@              �?               @               @       @                       @              �?333333D@�����ʜ@      �?              �?             �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333s9@fffff
�@                      �?      �?     �K@      �?              �?                                                       @      �?      �?33333CQ@33333�@      �?              �?      �?      R@              �?               @       @       @       @                       @              �?     �F@�������@      �?      �?      �?             �M@      �?              �?       @       @       @                              �?      �?      �?����̼T@ffff&'�@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@�����b@              �?                      @      �?                       @                                                      �?       @�����H@�����Eu@      �?              �?      �?     @P@      �?       @      �?                       @       @       @       @       @      �?        fffffZ@����,�@                      �?      �?      @      �?              �?                                       @                      �?       @fffff6T@�����Av@      �?                              8@      �?       @      �?               @                       @                      �?      �?33333�V@����ա@      �?                             �P@      �?       @      �?       @       @       @       @       @       @      �?      �?        fffff�]@ffff&|�@      �?              �?      �?      O@      �?              �?       @       @       @       @       @       @       @              @�����	[@ffff���@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      �?33333�3@�����1`@      �?                              8@      �?       @      �?               @       @                                      �?        fffff6U@������@      �?                              �?      �?              �?                                                              �?      @fffff�Q@fffff�Q@                                     �G@      �?       @      �?               @       @               @       @              �?       @fffff�Z@�����@                                       @      �?              �?                                                                       @�����<Q@     �]@                                      :@      �?       @      �?                       @               @       @              �?              Y@ffff�O�@                              �?      .@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@������p@      �?                              @@      �?       @      �?               @                                              �?        fffffT@����LH�@      �?                              @@      �?       @      �?       @                       @                                        ������U@����̜�@      �?                              (@      �?              �?                       @               @       @      �?               @������W@     ��@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      �?ffffff3@ffffff3@                      �?      �?      R@      �?       @      �?       @       @       @               @       @       @              �?�����l[@����L��@      �?                              �?      �?                                                                                      @������F@������F@                      �?      �?      @              �?                                                                      �?       @33333�8@������b@      �?                             �I@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333s4@�����J�@              �?      �?              <@      �?       @      �?                               @       @       @              �?      �?33333SY@fffff��@                      �?      �?      .@      �?                                                                                       @fffff&G@�������@      �?      �?      �?              4@      �?              �?               @                                              �?       @�����iR@     ޖ@      �?      �?      �?               @      �?              �?                       @                                      �?       @����̌R@33333�a@              �?                      @      �?       @      �?               @                       @       @              �?       @     �X@����̄�@      �?                              F@      �?               @      �?      �?      �?      �?      �?      �?       @              �?ffffff4@fffffL�@      �?      �?      �?      �?      @@      �?              �?               @                       @       @              �?      @�����|W@ffff�Z�@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @33333s3@33333s3@      �?              �?      �?     �P@      �?                       @       @       @       @                       @              @fffffvP@�����@                      �?              <@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @����̌9@������@      �?                              �?      �?                                                                              �?       @33333�F@33333�F@      �?              �?      �?     �F@      �?       @      �?               @       @                       @              �?        ������W@ffff�h�@      �?                              :@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ������3@�����}}@      �?                              D@              �?               @       @       @               @       @      �?              �?fffffO@������@      �?      �?      �?              P@      �?              �?       @               @                              �?              �?33333T@3333���@                                     �P@      �?               @      �?      �?      �?      �?      �?      �?      �?               @����̌4@�������@                      �?             �Q@              �?               @       @       @       @       @       @      �?                33333�P@ffff&Q�@      �?      �?      �?             �Q@      �?              �?               @       @       @               @       @      �?      �?     �W@ffff&3�@                                       @      �?              �?       @       @               @                              �?       @     �U@����̴f@      �?      �?      �?              O@      �?       @      �?               @       @               @       @      �?      �?       @     �Y@����Y�@              �?      �?      �?      <@              �?                       @                               @      �?      �?       @����̌C@fffff"�@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@������L@                                      6@      �?       @      �?                                       @                      �?        �����	U@�����w�@                      �?      �?     �M@      �?       @                               @       @       @               @      �?        fffffR@�����b�@                      �?      �?      R@      �?       @               @       @               @                       @              �?     �P@����L��@                      �?              .@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @3333339@fffff>x@      �?              �?             �C@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        33333s4@     ��@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y4@�����Y4@      �?                              @      �?              �?                       @                                      �?       @�����yR@������q@      �?              �?      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?33333�9@33333ʚ@                                      �?      �?                                                                              �?      @33333�F@33333�F@      �?              �?      �?     �O@              �?                       @       @       @                       @                ����̬C@������@      �?                              �?      �?                                                                                       @fffff�F@fffff�F@                      �?      �?     �P@      �?       @      �?               @               @       @               @              �?fffff�W@����̞�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @     @4@     @4@                      �?      �?     �D@      �?       @      �?               @       @       @       @       @      �?      �?        fffffF[@    @f�@                      �?             �L@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�3@fffffn�@      �?              �?      �?      I@              �?               @                               @                      �?      �?������C@fffff��@      �?                              @      �?              �?               @                               @                       @33333U@�����am@                              �?      <@      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@����̺�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                       @������2@������2@                      �?              @      �?                                                                                      @33333�F@333337t@      �?              �?               @      �?              �?       @                                                      �?      @     �R@����̐�@      �?              �?      �?      @      �?                       @               @       @               @              �?      �?fffff�Q@     �@              �?                      @      �?              �?                                               @                       @����̼S@fffff�w@      �?                              H@      �?               @      �?      �?      �?      �?      �?      �?      �?                33333�3@     d�@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?                      �?fffff�3@     8e@      �?              �?      �?      I@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @33333�8@����̵�@                                     �N@              �?               @       @       @       @                      �?              �?������E@�����@      �?              �?      �?      J@      �?       @      �?               @               @               @              �?             PW@3333��@      �?              �?              I@      �?       @      �?       @               @               @       @      �?      �?       @������Y@����Lo�@      �?                      �?      7@              �?               @               @       @                       @              @�����D@     Ί@                                     �B@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @������3@fffff��@      �?              �?      �?      :@      �?       @      �?                                       @                      �?       @     �T@33333-�@      �?                              ;@      �?                       @                       @                                      @������J@�����Ֆ@      �?              �?             �Q@      �?       @      �?               @       @               @              �?      �?             �W@ffff�ʹ@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @����̌3@����̌3@      �?                              ;@      �?               @      �?      �?      �?      �?      �?      �?              �?       @ffffff3@fffff��@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?       @                     �4@�����[�@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?33333�\@������@      �?              �?             �P@      �?       @      �?               @       @               @       @              �?      �?     @Z@    @ݻ@                                      �?      �?                               @                                                       @fffffFI@fffffFI@                      �?              R@      �?       @      �?       @       @       @               @       @       @      �?       @33333c[@�����@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @      �?      �?fffff�V@�����)�@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?                       @fffff&4@������V@                                      �?      �?                                                                              �?        33333sF@33333sF@                      �?              5@      �?       @      �?       @               @               @       @              �?        �����Z@    �0�@      �?              �?      �?      *@      �?              �?                       @               @       @              �?      @�����)X@fffff+�@      �?                              5@      �?       @      �?               @                                              �?       @fffff�T@fffff�@                      �?      �?      A@      �?                       @       @       @                              �?      �?      @ffffffN@33333�@      �?              �?              .@      �?       @      �?                       @               @       @              �?       @fffffFY@33333��@                                       @      �?       @      �?                       @               @       @              �?       @������X@     ��@                                      &@      �?       @      �?                                                                       @     �R@33333ŋ@                                      �?      �?              �?                       @               @                      �?       @�����\U@�����\U@      �?      �?      �?              R@      �?              �?       @       @               @                       @      �?      �?333333U@ffff���@                      �?      �?     �K@      �?       @               @       @               @               @      �?      �?             �R@    @��@      �?                             @Q@      �?       @               @       @       @       @               @       @      �?      �?     `T@    @��@                      �?             �E@      �?       @      �?       @       @                               @              �?       @fffff�W@����L�@      �?      �?      �?             @Q@      �?       @      �?               @                       @                      �?       @�����|V@ffff&��@                      �?              M@      �?       @      �?               @       @                       @      �?      �?       @33333�W@ffff&�@                                      @      �?              �?               @       @       @       @       @      �?      �?       @�����iZ@fffff�{@      �?              �?      �?      O@      �?       @      �?       @       @                       @              �?      �?      �?����̼W@����ٟ�@      �?                              M@      �?       @      �?                               @                                        �����)T@����Yǲ@      �?                              4@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?������3@fffffBv@      �?              �?              R@      �?       @               @       @       @       @       @       @       @      �?      �?      W@ffff&~�@      �?      �?      �?              L@      �?                       @       @       @       @       @       @       @      �?        �����iU@3333sز@                      �?              D@      �?       @                       @                                                      �?�����LL@33333��@                                      ;@      �?                               @               @                              �?      @33333L@fffff}�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�3@ffffffC@      �?              �?      �?     �E@              �?                       @                                                      �?�����L=@33333 �@                      �?      �?      I@      �?       @               @       @       @       @               @      �?      �?        33333T@fffff��@      �?                      �?      R@              �?               @       @       @       @       @       @       @              �?������P@3333�?�@      �?                              @              �?                                                                              @�����L8@�����Y@      �?                              1@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        fffff�3@������u@      �?                              4@      �?                                               @                                      @      I@fffffX�@      �?      �?      �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@����̱�@                      �?             �K@      �?       @               @       @               @                      �?      �?      �?33333�P@33333�@      �?              �?             �B@      �?       @               @                                                      �?      @fffff�K@     ��@      �?              �?             �Q@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff]@ffffF;�@      �?      �?      �?              D@      �?                                                               @      �?               @fffff�K@�����֡@      �?                              (@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?33333�8@fffff�q@                      �?              .@      �?               @      �?      �?      �?      �?      �?      �?                      �?33333s4@����̬t@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?33333�4@     �T@                                      �?      �?                                                               @              �?       @33333�K@33333�K@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?333333]@    `��@      �?                              .@      �?       @      �?               @               @               @                       @������W@fffff��@                                      @              �?                       @                               @              �?      �?�����D@�����Tr@                      �?      �?     �N@              �?                       @       @       @       @               @              �?����̬I@�����X�@              �?      �?      �?      D@      �?       @      �?                                       @       @              �?      �?33333�W@ffff�p�@      �?                             �A@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                333333:@33333׍@      �?                              &@      �?              �?                                                                       @����̌Q@fffff��@      �?                              @      �?              �?               @       @       @       @       @              �?       @������Z@������s@      �?              �?      �?     �F@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @33333s8@     �@      �?              �?      �?      ;@              �?                       @       @                       @      �?      �?      �?������F@�����y�@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@������3@                      �?      �?      R@      �?       @      �?       @       @       @       @               @       @              �?������Z@����L�@      �?              �?              J@      �?       @      �?       @               @       @                       @      �?      �?fffff�V@������@                                      =@      �?       @      �?                       @               @       @              �?      �?fffff�X@fffff�@      �?                              *@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����L3@fffff:p@                      �?              *@              �?                               @               @       @              �?             `H@33333˃@                      �?      �?     �I@      �?                       @       @       @       @       @       @       @              �?     `U@3333�E�@              �?                      G@      �?       @      �?               @       @               @       @              �?       @�����Z@�������@                      �?             �H@      �?              �?               @       @               @       @                       @������X@     ��@                                      ,@      �?                               @                                                       @�����9I@������@                      �?              P@      �?                               @       @       @               @       @      �?      @33333Q@������@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      �?�����Y4@����̌A@      �?                               @      �?       @      �?       @                                       @                      @     �V@     �e@                      �?      �?     �K@      �?       @               @       @               @       @              �?      �?      �?     �R@ffff�u�@      �?              �?      �?      M@      �?       @               @       @       @       @                       @              �?fffff�Q@    @��@      �?      �?      �?              @              �?                               @                                      �?       @fffff�=@     �]@      �?                              1@      �?       @      �?                       @       @                      �?               @     �U@     	�@      �?                      �?      ,@      �?                       @       @       @       @               @       @                fffffS@33333{�@      �?                              K@      �?                       @       @                       @               @      �?        33333SP@�����q�@      �?      �?                      @      �?       @      �?               @                               @              �?       @33333sV@�����i@      �?              �?             �E@      �?                                                       @              �?      �?      @�����,L@����L��@      �?              �?              &@      �?                                                                              �?        33333�F@33333O�@                                      �?      �?              �?                                                              �?      @����̬Q@����̬Q@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����5@�����5@      �?                              �?      �?       @                               @                                               @�����,K@�����,K@      �?              �?              &@      �?       @      �?                                                              �?       @����̼R@�����͉@              �?                      @      �?       @      �?                                       @                      �?      �?������T@������{@      �?                              �?      �?                                                                                      @fffff&G@fffff&G@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@33333s[@      �?              �?      �?      �?      �?              �?                                               @              �?       @33333CT@33333CT@                      �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�3@33333Օ@      �?              �?              $@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������3@fffff�g@                                      .@      �?       @               @                                       @              �?        �����)P@fffff�@                                       @      �?                       @                       @               @                        33333�P@     �@              �?                      R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?fffffV]@     z�@      �?              �?      �?      Q@      �?       @      �?       @       @       @       @       @       @       @      �?        ����̬\@����٩�@      �?      �?      �?              @@      �?       @      �?                                                              �?       @������R@3333���@      �?                              K@      �?              �?       @               @       @                      �?               @�����U@������@      �?      �?                     �P@      �?              �?       @       @               @       @       @       @      �?       @33333CZ@3333��@                      �?      �?     �O@      �?                       @                                               @      �?        33333SI@    �*�@      �?              �?      �?     @P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     �8@fffff̚@      �?              �?              R@      �?       @      �?               @       @               @       @       @      �?        33333�Z@����Y��@      �?                              (@      �?       @      �?               @       @       @       @       @              �?      @�����<\@     ��@      �?      �?      �?             �F@      �?       @      �?               @       @       @       @              �?      �?        ����̬X@����̭�@      �?      �?                      "@      �?       @      �?                       @               @       @              �?       @      Y@����̴�@                                      �?      �?                                       @       @       @       @      �?              �?fffff�R@fffff�R@                                      N@      �?       @               @               @       @                      �?               @     0P@     ��@      �?                              2@      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@     hv@      �?      �?      �?              @      �?       @      �?                       @               @       @              �?       @�����|Y@������@      �?                              6@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@     hz@                      �?      �?     �P@      �?       @      �?                       @       @       @       @       @      �?        �����iZ@ffff�=�@      �?                              J@      �?              �?                       @                       @              �?      �?33333�T@fffff�@      �?                              >@      �?              �?                                       @       @              �?       @     �V@3333���@                      �?      �?      Q@              �?                       @       @       @       @       @       @              �?fffff&N@     �@              �?                      K@      �?       @                       @               @       @              �?              @fffffR@����\�@                      �?      �?      "@      �?              �?                               @                              �?       @fffff�R@     <�@      �?                              I@      �?       @                               @       @               @       @                     `Q@fffff��@      �?      �?      �?             �N@      �?       @      �?               @               @                      �?      �?        33333cU@    ���@      �?              �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        3333339@������@      �?      �?      �?              M@      �?       @      �?       @       @       @               @       @      �?      �?       @fffff6[@    @��@      �?                             �C@      �?              �?                       @       @                      �?               @�����yT@    �'�@      �?              �?      �?      A@      �?               @      �?      �?      �?      �?      �?      �?                      @������4@33333߃@      �?              �?      �?      D@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@�����G�@                      �?      �?      R@      �?       @               @       @       @       @       @       @       @              �?����̼V@3333s��@      �?                              @      �?                                                                                      @fffffFF@     �k@      �?                              �?      �?              �?                                       @       @              �?       @33333�V@33333�V@                      �?      �?      R@              �?                       @               @       @       @       @              �?33333�J@     ��@                                      =@              �?               @       @               @                      �?              �?     �C@     �@      �?                              4@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�3@fffff6z@      �?              �?      �?      *@      �?              �?                       @               @       @                       @     @X@�����ٔ@      �?              �?             �I@      �?                       @       @       @       @       @       @       @      �?      �?     �T@ffff��@      �?      �?      �?              ?@      �?       @      �?       @                               @                               @�����\V@����L�@      �?              �?      �?      Q@      �?                       @       @               @       @       @       @                fffff�T@3333s��@      �?              �?             �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������8@     ��@                                      .@      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?ffffff9@������x@                      �?      �?      R@      �?       @               @       @       @               @       @       @      �?      �?fffff�T@����LG�@      �?                              O@      �?       @               @       @       @       @                       @                �����YQ@    ���@      �?                              $@      �?       @               @                                                      �?      �?     @K@�������@      �?              �?              R@              �?               @       @       @                               @                �����E@     $�@                                     �N@      �?       @                       @       @       @       @       @       @              �?�����)V@    @ɴ@      �?                              �?      �?              �?                               @                                       @     �R@     �R@      �?              �?      �?      �?      �?              �?                                                              �?       @     �Q@     �Q@      �?              �?      �?     �F@      �?       @               @       @               @       @               @              �?fffffvR@     V�@      �?              �?      �?      �?      �?              �?               @                                                      �?fffff�R@fffff�R@              �?                     �A@      �?       @      �?       @                               @       @              �?       @33333�X@33333ū@      �?                              @      �?                               @                       @                               @������M@�����Yv@                      �?      �?     �L@      �?              �?               @                       @       @      �?      �?       @     �W@����̟�@                                      @      �?              �?                                       @                      �?      �?     @T@�����Yx@                      �?             �M@      �?              �?       @               @                              �?      �?      �?     PT@3333s�@              �?                     �K@      �?       @      �?                       @               @       @      �?      �?       @�����	Y@    �!�@                                     �A@      �?               @      �?      �?      �?      �?      �?      �?                             @3@33333M�@                                      <@      �?              �?                                               @              �?       @fffff&T@ffff扡@                      �?      �?     @P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����L9@33333R�@      �?                              7@      �?       @      �?                       @       @       @                      �?      �?�����9X@ffff�J�@      �?                              @      �?              �?                       @                       @                      �?�����lU@     p@      �?              �?      �?       @      �?                                                                              �?       @     @F@33333�V@      �?      �?      �?              F@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�����Y3@     z�@                                      7@      �?       @      �?               @                       @       @              �?      �?����̬X@33333��@                      �?      �?     @P@      �?       @                       @               @       @       @       @      �?        ������S@ffff�ϳ@                      �?      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@33333�@                                      @      �?                                               @       @                      �?      @     �M@33333�y@                      �?      �?      P@      �?       @               @       @       @       @       @       @       @      �?      @fffff�V@3333s��@      �?              �?      �?      1@      �?              �?                                                              �?       @     @Q@�������@                      �?              (@      �?                               @                                              �?       @     �I@����� �@                                      @      �?       @      �?                                       @       @              �?        33333cW@33333À@                      �?              �?      �?                                                                              �?       @     �F@     �F@      �?                              $@      �?                       @                       @       @                                      O@�����'�@      �?              �?             �I@      �?       @                                       @       @       @       @      �?        ������R@    �z�@                      �?      �?     @Q@      �?       @      �?               @       @               @       @              �?       @������Y@ffff��@      �?                      �?      >@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �����Y9@fffff��@      �?              �?              E@      �?               @      �?      �?      �?      �?      �?      �?       @               @     @4@     �@                                      ?@      �?       @      �?                       @                       @              �?       @�����yV@������@                                      E@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @fffff�4@�������@      �?                              �?      �?                                                                              �?        fffffF@fffffF@      �?              �?              L@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?33333�3@     ��@                      �?      �?      A@      �?                       @       @       @       @       @       @       @              @     0U@ffff�.�@                                      @      �?                                       @               @       @      �?      �?       @�����|Q@fffff�k@                                       @      �?       @      �?                                       @       @              �?       @������W@����̜h@      �?              �?              2@      �?       @      �?                                       @       @              �?       @����̬W@�����_�@      �?                              @@      �?                                                       @       @      �?      �?        fffff6P@�����k�@                      �?      �?     �O@      �?                       @       @       @       @                       @              @fffff�O@fffff\�@                      �?      �?     �G@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����4@�����ŏ@                      �?      �?      $@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff&4@������k@      �?              �?              @      �?       @      �?                                                              �?       @     �R@     `{@      �?                      �?      8@              �?               @                       @                       @              @     �A@fffff��@                      �?      �?      P@      �?       @      �?       @                       @       @       @      �?      �?        �����Z@�����A�@                      �?      �?      6@      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@�����y@                      �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@������q@      �?              �?      �?      J@      �?                               @       @       @       @              �?      �?       @     0Q@3333�5�@      �?      �?                     �P@      �?       @      �?               @       @       @       @       @      �?              �?������[@�����@                      �?      �?      H@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�4@     ��@      �?                              3@      �?              �?                               @               @      �?      �?      �?������U@�������@                                     �C@      �?                                               @               @      �?               @fffff�M@����LB�@              �?                      7@      �?              �?       @                                                      �?        ������R@33333��@              �?      �?             �C@      �?       @      �?                               @       @       @              �?       @     PY@����Lڮ@      �?              �?              8@      �?       @      �?                       @               @       @              �?       @33333CY@�������@                                      @      �?       @      �?                       @       @                              �?       @     �T@     z@                                       @      �?                       @                               @                      �?       @      N@     |~@                                      <@      �?       @      �?               @                               @              �?       @�����|V@������@      �?              �?              �?      �?              �?                                                              �?       @�����IQ@�����IQ@      �?              �?      �?     �N@      �?               @      �?      �?      �?      �?      �?      �?      �?              @ffffff4@�����)�@      �?                              (@      �?       @      �?                                       @       @              �?       @33333X@fffff�@                      �?              F@      �?                       @       @       @                              �?      �?      @     �N@fffffD�@                                      J@      �?       @               @               @       @       @              �?              �?     �R@����LK�@                      �?      �?      �?      �?              �?               @                                              �?       @����̬R@����̬R@      �?              �?              R@      �?       @      �?       @       @       @       @               @       @                ffffffZ@    ���@      �?              �?             �I@              �?                       @                                              �?      �?�����>@������@              �?      �?             �P@      �?       @      �?                       @       @       @       @      �?      �?      �?�����|Z@    @?�@      �?                              �?      �?       @      �?                                       @                               @      U@      U@              �?      �?              :@      �?              �?                       @               @                      �?      �?�����lU@     &�@      �?                              >@      �?                       @               @                               @      �?      @33333�K@fffffי@      �?              �?      �?      I@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�����Y4@�����W�@      �?                              $@      �?              �?       @               @               @       @      �?      �?       @������X@����̣�@                                     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?      �?������[@3333�s�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                        �����4@�����4@                      �?      �?      @      �?       @                                                                               @ffffffH@������u@      �?                              M@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        fffff&3@     .�@      �?                              L@      �?       @      �?               @               @               @              �?       @����̜W@������@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@     H`@                                      ;@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������3@33333��@      �?                              �?      �?       @      �?                                                              �?       @������R@������R@                      �?              3@      �?       @      �?                                       @                      �?       @fffff�U@�����q�@                      �?      �?     �P@      �?       @      �?       @                       @               @      �?      �?      �?fffff�W@3333sŸ@                                       @      �?               @      �?      �?      �?      �?      �?      �?                       @fffff�3@33333�L@      �?              �?      �?      1@      �?       @               @                       @                      �?      �?      @�����O@�����"�@                                      (@      �?       @      �?                       @               @       @              �?        �����	Y@333331�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @33333s4@33333s4@      �?                              H@      �?       @      �?               @       @               @       @       @      �?        fffff[@3333s˳@                                     �O@      �?              �?                       @       @       @              �?      �?      �?33333�V@     ��@                                     �K@      �?                       @                                                      �?      �?fffffFI@    �!�@      �?                               @      �?                                                                                      @fffff�E@fffff�t@              �?      �?              &@      �?       @      �?                       @       @       @       @              �?        33333Z@�������@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @������4@33333sO@      �?                              8@      �?                               @                                              �?      @������H@     	�@                                      >@      �?              �?                               @       @       @      �?      �?        ������W@33333��@      �?                              @      �?              �?                                                                        �����IQ@fffff�~@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@fffffY@              �?      �?              5@      �?       @                       @       @                       @      �?                ������Q@33333d�@                      �?      �?     �I@      �?       @      �?       @       @                               @              �?       @33333sW@����Y��@      �?                             �J@              �?               @       @                               @              �?        fffff&G@3333��@                      �?      �?     �E@      �?                               @                                                      @�����I@������@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                        fffff�3@fffff�3@                                      2@      �?       @                                                                      �?       @fffff&I@fffff��@                      �?      �?      A@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?33333�8@fffff�@                      �?      �?      J@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@33333��@                      �?      �?     �P@              �?               @       @                                       @                33333B@ffff��@                      �?      �?      @      �?                       @                                                              @�����YI@������u@      �?                      �?     �N@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@����̐�@      �?              �?      �?      F@              �?               @       @       @       @               @       @      �?      �?fffffK@fffff��@              �?      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?        ������\@�����F�@      �?      �?                      @      �?       @      �?                                       @                      �?       @333333U@������@                      �?             �Q@      �?       @      �?               @       @               @       @       @      �?        �����IZ@     ��@      �?              �?             �P@              �?               @       @       @       @       @               @      �?        �����LL@fffff��@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?                      �?     �3@fffffnr@                                      (@      �?       @      �?                               @                              �?      �?33333�S@     �@                                      6@      �?       @      �?                               @       @                      �?       @     �V@33333'�@                                      @      �?              �?                                       @                      �?       @������S@fffffP�@              �?      �?             �P@      �?       @      �?       @       @                       @       @      �?      �?       @ffffffZ@ffff&Ȼ@      �?                              @      �?                               @                                              �?      @33333�H@33333C`@                                      @      �?       @      �?                                                              �?       @������R@������r@                      �?      �?      R@      �?       @               @               @       @       @       @       @      �?      �?�����yU@    �޷@      �?              �?      �?     @Q@      �?              �?               @               @       @               @      �?      @�����	W@ffff�P�@      �?      �?      �?             �B@      �?              �?                                                              �?             R@ffff��@      �?              �?              �?              �?                               @               @       @              �?       @�����,I@�����,I@                                      @      �?              �?                                                              �?      @�����yQ@�����@                      �?              I@      �?       @                               @               @       @      �?                ������R@fffffH�@      �?              �?      �?      K@      �?       @               @       @               @                       @      �?      �?�����iP@fffffݫ@              �?                       @      �?              �?                                               @              �?       @fffff�S@�����ah@      �?                      �?      L@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @3333335@�����Z�@      �?      �?                     �D@      �?       @      �?                       @               @       @              �?       @������X@    �[�@                                     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�����:@33333~�@      �?                             �F@      �?                       @               @               @       @              �?       @������R@�������@      �?                      �?     �G@      �?                       @       @                                              �?       @fffff�K@������@      �?              �?      �?      6@      �?               @      �?      �?      �?      �?      �?      �?      �?                     @4@     �~@      �?                              <@      �?       @      �?       @       @                               @              �?      �?     �W@�����Ƥ@      �?                             �A@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @������9@     *�@      �?                      �?      3@              �?                                                                      �?      �?�����Y9@����̰�@                              �?      @      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @33333s9@�����U@      �?              �?             �H@              �?                       @                       @       @       @              �?33333�H@�����Ӣ@              �?      �?             �J@      �?              �?               @       @       @       @              �?      �?       @     �W@3333s�@      �?              �?      �?     �Q@      �?                       @               @       @               @       @      �?      �?fffff�Q@fffffm�@      �?              �?      �?      R@      �?                       @       @               @       @               @                �����Q@����Y��@      �?                              @      �?                                       @                                      �?       @33333�H@�����!e@      �?              �?             �P@      �?       @               @       @       @                               @      �?      �?fffff�P@3333sL�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @������4@������4@      �?      �?      �?              @      �?       @      �?                       @                                      �?       @333333T@������|@                                       @      �?              �?                                       @                      �?       @     �S@     �d@              �?                      ,@      �?       @      �?               @                                              �?       @����̼S@fffff7�@      �?      �?                      @      �?              �?                                       @       @              �?       @     `V@33333�}@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@fffff��@      �?              �?             �N@      �?       @      �?               @       @       @       @       @              �?       @fffff�\@ffff&ܻ@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        �����L7@�����\�@              �?      �?             �K@      �?       @      �?               @       @       @                                       @����̜V@����̴�@                      �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @3333334@fffffP�@      �?              �?      �?      G@      �?       @      �?               @                                              �?              T@fffffs�@                      �?              8@      �?       @      �?                                                              �?      �?������R@fffffO�@                                      �?      �?       @      �?                                               @              �?       @     @U@     @U@              �?      �?             @P@      �?              �?               @       @       @       @       @       @      �?      �?fffffvZ@    �E�@                      �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @                fffff�\@    @��@      �?              �?              ?@      �?       @      �?                       @               @                              �?�����)V@fffff��@              �?                      0@      �?                                               @       @                               @33333�M@33333��@                      �?              M@      �?       @      �?       @       @       @               @       @       @      �?        �����\[@���̌ �@                      �?      �?      J@      �?              �?       @               @       @                              �?        33333U@������@      �?                              O@              �?               @       @       @       @                       @      �?        ������E@�����t�@                                      "@      �?       @      �?                                                              �?      �?������R@�����΃@                      �?      �?      @@      �?       @      �?               @                       @       @              �?       @fffff�X@33333#�@                      �?               @              �?                                                       @              �?       @����̌A@     0Q@      �?                              �?      �?              �?                                                              �?       @�����yQ@�����yQ@                                       @      �?       @      �?                                       @                      �?       @33333�U@�����Ї@                      �?      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @     �3@      q@              �?                      5@      �?       @      �?                                       @       @              �?        ������W@fffff��@                      �?              "@      �?              �?                                       @       @                       @�����\V@����̨�@                      �?      �?      7@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����9@������@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?fffff�3@33333W@      �?                              :@      �?               @      �?      �?      �?      �?      �?      �?      �?              @ffffff3@fffffl�@      �?      �?                     �@@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        fffff�8@fffff~�@              �?      �?              (@      �?       @      �?               @       @               @                      �?       @fffff�X@����̐�@      �?      �?                      *@      �?                               @                       @                      �?       @33333�M@����̢�@                      �?      �?       @      �?              �?               @                                              �?        33333cR@�����,b@      �?                               @      �?              �?                       @               @       @                       @����̼W@33333Cf@              �?                      @      �?              �?       @                                                                �����S@�����y@      �?                              @      �?              �?                               @       @       @              �?       @fffffX@fffffV|@      �?              �?      �?     �C@      �?       @      �?                       @               @       @      �?               @      Y@������@                      �?             @Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     @8@33333��@      �?              �?             �A@              �?               @               @               @       @      �?              �?33333�J@�����+�@                                      :@              �?                               @       @       @                      �?      �?�����9F@33333�@      �?              �?      �?      @@              �?                               @               @       @                      �?�����LI@�����ՙ@                                      �?      �?              �?       @       @               @                              �?      @������T@������T@      �?                              5@              �?                       @               @                              �?      @      B@33333a�@                                      <@              �?                               @       @                              �?      @     �A@33333�@                      �?      �?      $@      �?                               @       @                                      �?      @fffff�K@fffff:�@              �?      �?              L@      �?       @               @       @       @       @                      �?      �?      �?�����Q@     \�@                              �?      @              �?               @       @       @               @       @              �?      @������L@     �k@      �?              �?              8@      �?       @      �?               @       @               @       @              �?       @�����)Z@ffff�ܣ@                      �?              8@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff&4@������|@              �?                      �?      �?              �?                                       @       @              �?       @33333�V@33333�V@                      �?               @      �?       @      �?                                       @                      �?       @33333U@������`@                      �?      �?     �@@      �?              �?                       @               @       @      �?      �?       @33333sW@     i�@                                       @      �?              �?                                                              �?       @����̬Q@������b@              �?                      �?      �?              �?                       @                       @              �?       @     @U@     @U@      �?                              F@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?     �3@     �@      �?                              L@      �?       @      �?               @                       @       @                       @fffff�X@����͵@                                     �A@      �?       @      �?                       @               @       @              �?       @     Y@33333��@                                       @      �?                       @                       @                      �?                      K@     �{@      �?                              K@              �?               @       @                               @       @                �����G@ffff���@                                      $@      �?               @      �?      �?      �?      �?      �?      �?                      @������2@ffffffd@      �?                      �?      J@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?fffff�3@33333�@      �?              �?      �?      ,@      �?                       @       @                       @                      �?       @�����\P@�����L�@      �?      �?      �?              $@      �?       @      �?                                               @                       @33333cU@     ��@      �?              �?              M@      �?                       @       @       @                              �?              �?fffff&N@�����׫@                      �?      �?     �P@      �?       @               @                               @       @       @      �?       @     �R@3333sm�@                                      @              �?                                       @       @       @      �?      �?      @     �H@33333�o@      �?              �?      �?     �C@      �?              �?               @                       @                      �?      @33333�U@     ��@                      �?      �?     �E@              �?               @               @       @       @       @      �?      �?      �?333333N@������@                                     �N@      �?       @      �?                       @                       @                      @�����LV@�����|�@              �?                     �F@      �?       @               @                       @               @              �?       @33333�Q@ffff��@      �?                              G@      �?                                                                              �?      �?������F@����L"�@              �?      �?              :@      �?       @      �?                       @               @       @              �?        fffff�X@fffff��@      �?              �?              L@              �?                               @       @       @       @      �?      �?        fffffK@������@      �?                             �D@      �?       @                               @                       @      �?              @     @P@�����ǣ@              �?                      @      �?              �?                                                              �?       @������Q@fffff�i@              �?      �?             �E@      �?       @      �?       @               @       @       @       @      �?      �?      @33333c[@    @޲@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                        3333334@�����LI@      �?                              @      �?                                       @       @       @       @                        ������R@fffff�x@      �?              �?             �Q@      �?       @      �?       @               @       @       @       @       @      �?      �?33333#[@     ��@      �?              �?      �?      R@      �?       @               @               @       @                       @      �?      �?     �P@�����˲@      �?              �?              N@      �?       @      �?                       @               @       @       @              �?�����IY@fffff��@                                      (@      �?                                                                              �?             �F@�����b�@      �?      �?                      �?      �?       @      �?                                                              �?       @�����S@�����S@      �?              �?      �?      Q@      �?       @               @       @       @       @       @       @       @      �?      �?�����W@�������@      �?                              @      �?       @      �?               @       @                       @                       @33333#X@�����A@                      �?      �?      4@      �?       @      �?                       @       @               @              �?             �W@������@                      �?              P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?      9@33333Ø@      �?              �?      �?      "@      �?                               @               @                                      @ffffffK@�����L|@      �?      �?      �?              @@      �?       @      �?                                               @                       @33333SU@33333ʤ@              �?      �?              F@      �?       @      �?                       @       @       @       @                       @�����	Z@ffff���@                      �?      �?     �K@      �?       @      �?       @       @                                              �?       @fffffFU@3333���@                              �?     �O@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �3@fffff��@      �?              �?      �?     �Q@      �?       @      �?       @               @               @       @       @               @33333cZ@    ��@      �?      �?      �?      �?      A@      �?       @      �?               @       @       @       @       @              �?       @�����9[@fffffR�@              �?                       @              �?                                                                               @�����Y8@������D@      �?                              =@      �?                                       @       @       @       @      �?      �?        fffff�R@����̇�@      �?                              8@      �?                       @                       @                                       @�����yK@     �@                                      2@      �?       @      �?                                       @                      �?       @�����LU@�����G�@              �?      �?      �?      A@      �?       @      �?               @                                              �?      @fffff�S@�����<�@      �?                              @      �?       @      �?                                       @       @                       @�����X@�������@                                      &@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����4@fffff�m@      �?              �?             �P@      �?       @      �?       @       @       @       @       @       @      �?                33333�\@ffff&�@                                     �D@      �?                       @               @       @       @       @      �?      �?        fffff�S@    ��@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        fffffF\@    @�@                      �?             �N@      �?       @      �?                               @       @       @      �?                �����IY@ffff��@                                      B@      �?       @      �?               @                       @       @              �?       @������X@33333?�@                      �?      �?      K@      �?       @                       @       @       @       @       @              �?       @����̌U@������@      �?                      �?      $@      �?       @      �?                                       @       @                       @������W@33333�@      �?      �?      �?             �K@      �?       @      �?                                                              �?       @     �R@����̨�@                                      @      �?              �?                       @       @               @              �?       @     PV@�����p~@      �?              �?              9@      �?       @                               @                                              �?fffff�K@33333��@      �?                              �?      �?              �?                                       @       @              �?       @fffffV@fffffV@      �?      �?                      C@      �?                               @       @       @       @              �?      �?      �?������Q@3333���@      �?              �?      �?       @      �?                       @       @               @                       @              @     �M@     P`@      �?                              �?      �?              �?                                               @              �?       @333333T@333333T@                                      >@      �?                       @                                                      �?      @ffffffH@     �@      �?      �?      �?             �E@      �?              �?               @       @               @       @      �?      �?        33333#Y@     а@      �?              �?              "@      �?              �?               @       @       @       @                      �?      @fffff�W@�����ԋ@      �?              �?      �?     @P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?������3@33333̓@                      �?              5@      �?       @      �?                                       @       @              �?       @33333�W@fffffq�@                                      @      �?                                                                              �?      @      G@333333h@      �?                              @      �?              �?       @                       @                              �?      @33333�T@������j@      �?              �?             �Q@      �?       @                       @       @       @       @               @              �?fffffS@    @��@                      �?      �?      <@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@     ��@      �?                              @      �?       @      �?                                                              �?       @33333S@fffff�s@                      �?      �?     �G@      �?       @               @       @               @       @       @       @      �?      �?33333SU@    @�@                              �?      1@      �?       @      �?               @       @       @                              �?      �?�����,W@fffffS�@      �?      �?      �?             �L@      �?       @      �?               @                               @              �?       @fffffvV@����Y=�@                      �?      �?      @              �?                       @               @                                       @      A@�����qd@      �?              �?              N@      �?              �?               @                       @       @      �?      �?       @������W@    @�@                      �?             �J@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����3@������@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?       @              @33333s3@33333�d@                                      1@      �?       @      �?                       @                                                33333T@������@                                      (@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        �����Y3@33333kk@                      �?               @      �?              �?               @       @                                                ������S@     �d@      �?              �?      �?      ;@      �?              �?       @       @                                      �?      �?      �?�����)T@    �C�@                      �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?                      @������3@33333q@                                     �B@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@     ��@                                      :@      �?              �?                                       @       @              �?        333333V@3333�ġ@      �?      �?      �?      �?      N@      �?       @      �?       @       @                               @              �?       @     PW@���̌��@                                      @      �?       @      �?               @                                              �?        33333�S@�����W�@                      �?      �?      G@              �?               @       @                                                        fffff�A@     Q�@                                       @      �?              �?                                                              �?       @������Q@33333�^@              �?                      L@      �?       @               @               @       @               @       @                     PR@fffff��@      �?      �?      �?              1@      �?       @      �?                                       @       @              �?       @33333�W@�����o�@      �?                              5@              �?               @                       @       @                      �?      @fffff�E@     ��@      �?              �?      �?      8@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����8@33333[�@                      �?      �?      O@      �?                       @               @       @       @              �?      �?             �Q@3333s��@      �?              �?             �Q@      �?              �?       @       @               @                       @                fffff&U@33333J�@      �?              �?      �?      4@      �?              �?                                                              �?       @����̜Q@�������@                                      &@      �?               @      �?      �?      �?      �?      �?      �?      �?              @      4@fffff~j@      �?              �?      �?      ,@      �?       @               @       @                               @                      @�����LQ@33333��@              �?      �?              1@      �?       @      �?       @               @                                      �?        fffffVU@�����ݖ@      �?              �?      �?      L@      �?       @      �?                       @       @       @       @       @      �?       @������Y@    ��@      �?              �?      �?      *@      �?                       @                                                      �?      @������H@�����[�@      �?                              $@      �?                               @                       @                      �?      @33333�M@�������@      �?                              "@      �?       @      �?               @                       @       @              �?      �?33333�X@     ��@                      �?              E@      �?       @       @      �?      �?      �?      �?      �?      �?       @               @     @9@�����P�@                                       @      �?       @                       @                                                      @33333K@�����iY@      �?              �?      �?     �F@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y4@�����	�@                                     �F@      �?       @      �?               @                       @                      �?      �?33333SV@3333�a�@      �?              �?             �Q@      �?       @      �?       @       @       @       @       @       @       @      �?       @     ]@    `��@      �?                             �L@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������2@fffff�@      �?      �?      �?             @Q@      �?       @      �?               @       @       @       @       @       @      �?        �����[@33333��@      �?                      �?      5@      �?                                                                                      @33333�F@fffffȎ@                                      .@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����4@33333�r@      �?                             �F@              �?               @               @       @                      �?                fffff&E@     Ü@                      �?      �?       @      �?                                                       @       @                      @�����lP@33333�`@      �?      �?      �?              @      �?       @      �?                       @               @       @              �?       @     �X@�����˄@      �?                              R@      �?       @      �?               @       @               @       @       @      �?        �����9Y@����#�@      �?                              �?              �?                                                                      �?       @     @8@     @8@                              �?     �P@      �?       @      �?               @               @       @       @      �?      �?        fffff�Z@3333�L�@      �?                              2@      �?               @      �?      �?      �?      �?      �?      �?                       @      3@������u@                                      M@      �?              �?       @       @       @               @       @      �?      �?       @����̜Z@������@      �?              �?             �@@      �?              �?                       @               @       @      �?      �?       @33333�W@    ���@      �?                              6@              �?                       @       @                       @      �?      �?             �E@�����<�@      �?              �?              1@      �?       @      �?               @                                              �?              T@������@      �?              �?              "@      �?                                       @               @       @              �?      @33333�Q@33333��@                                      &@      �?       @      �?                       @               @       @              �?        fffffvX@�����E�@      �?                      �?      9@              �?               @                               @              �?      �?      �?33333SD@fffffT�@                      �?      �?      E@      �?              �?                       @       @       @       @       @      �?       @�����Y@ffff�ϰ@      �?                              $@      �?              �?                       @               @       @              �?       @������W@fffffc�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                       @�����L3@�����L3@      �?              �?              2@      �?              �?                       @       @                                       @����̌S@     �@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @      �?      @�����YV@���̌�@                      �?             �N@      �?       @      �?                       @       @       @       @              �?       @fffff�Z@����Y_�@      �?                              *@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333s3@33333�p@      �?              �?      �?     �G@      �?       @                       @                                                       @      K@fffffԣ@      �?                              �?      �?                                       @                                      �?       @     @I@     @I@              �?                      5@              �?               @                               @                      �?       @33333�D@�����@�@      �?      �?                      @      �?       @      �?                                                              �?       @33333S@������l@      �?      �?      �?              *@      �?       @      �?       @       @                               @                      �?33333sW@     ��@      �?              �?             �J@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�3@33333X�@      �?                              @      �?       @      �?                                                              �?        �����R@�����s@              �?                     �A@              �?                               @               @                      �?       @������C@fffffj�@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?      �?                     �4@33333�S@      �?              �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                      9@�����+�@                      �?      �?      R@      �?       @      �?       @       @       @               @       @       @              �?33333c[@    @Ͼ@      �?      �?      �?             �P@      �?       @      �?               @               @       @       @       @                ������Y@3333�M�@              �?              �?      �?      �?              �?                                                              �?       @     �Q@     �Q@      �?                              &@      �?       @       @      �?      �?      �?      �?      �?      �?                      �?fffff&7@fffff�n@      �?                               @      �?              �?                       @               @       @              �?       @����̬W@fffff"�@      �?                      �?      7@      �?                               @               @                              �?        fffff�K@������@      �?      �?      �?              N@      �?       @      �?               @       @               @       @      �?      �?       @fffffZ@3333sø@      �?              �?             �Q@      �?       @                       @       @       @       @               @                �����<R@���̌��@      �?              �?      �?      &@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@     8l@                                      2@      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@33333{x@                              �?      I@      �?                       @               @       @       @              �?      �?      �?33333�Q@����L,�@      �?                      �?       @              �?               @                       @               @       @      �?      @fffffFF@33333wu@                                      ,@      �?       @      �?                       @                                      �?       @�����T@     ��@      �?                              E@      �?       @      �?       @       @       @                       @      �?      �?       @     �X@3333sʰ@                                      7@      �?                               @       @                              �?                fffff�K@fffff��@      �?                      �?      �?              �?                       @               @                                      @������@@������@@                      �?      �?     �E@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        33333s8@33333	�@              �?      �?             �P@              �?                       @       @               @              �?                fffff�F@    ���@              �?      �?             @P@      �?              �?       @       @       @                       @                       @������W@ffff&�@      �?                              L@      �?                               @               @       @       @      �?      �?             �R@ffff���@      �?              �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @                �����L4@������@      �?              �?      �?     �F@      �?       @      �?               @       @       @       @       @       @      �?             p[@ffff�$�@      �?              �?      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����L:@�����c�@      �?              �?      �?      L@              �?                       @       @                              �?      �?      �?�����B@     Ξ@                      �?              Q@      �?       @      �?       @       @       @       @       @       @       @              @fffff�]@����6�@              �?                      �?      �?       @      �?                                               @              �?       @33333CU@33333CU@                                      R@      �?       @      �?               @       @       @       @       @       @      �?      �?33333[@�����~�@              �?      �?              ;@      �?       @      �?       @                       @       @       @              �?        33333Z@    �g�@                                      �?              �?                                                              �?              @������9@������9@      �?                              �?      �?              �?                                                              �?       @33333sQ@33333sQ@      �?      �?      �?             �E@      �?       @      �?               @       @               @       @              �?       @     �Y@����L>�@                                       @      �?                                       @                       @                       @�����lN@������[@                      �?              G@      �?       @      �?               @               @       @       @      �?      �?       @������Y@ffff��@      �?              �?      �?      (@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@�����%p@      �?              �?      �?      >@      �?       @      �?               @               @                              �?        33333�T@fffff�@      �?      �?                      �?      �?       @      �?                                                              �?       @fffff�R@fffff�R@                                     �D@      �?       @               @               @       @               @              �?        ������R@����L%�@                                       @      �?              �?                                                              �?       @����̼Q@fffff>a@              �?      �?      �?      G@      �?       @      �?       @       @               @       @       @              �?       @����̌[@����l�@      �?      �?      �?              5@      �?                       @       @                               @              �?        �����<P@33333�@      �?      �?                      @      �?                                       @                                               @�����,I@     �m@                                      $@              �?               @                                                              @     �=@fffff�r@      �?                      �?      ;@      �?               @      �?      �?      �?      �?      �?      �?       @              @������4@�����.�@                                       @      �?                                       @       @               @                      @fffffP@����̀@                      �?              (@      �?       @               @               @               @       @      �?               @fffff�S@     f�@      �?              �?      �?      R@      �?       @      �?               @       @               @       @      �?      �?      �?�����Z@     #�@      �?              �?              I@      �?       @      �?               @                       @       @      �?      �?       @     �X@3333���@                      �?      �?      7@      �?       @      �?                                       @                      �?       @     �T@������@      �?              �?              .@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?33333s3@�����Mu@      �?      �?                      �?      �?                                                                              �?      @������F@������F@      �?      �?      �?             �P@      �?       @      �?       @       @                                                        fffff�T@�����Ե@      �?                              �?      �?                                                                                      �?�����G@�����G@                      �?              1@              �?                       @       @                                      �?      �?33333�A@fffff0�@      �?              �?             �Q@      �?                       @       @       @       @                       @              �?�����<P@    @��@      �?              �?      �?      5@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@������u@      �?              �?      �?      B@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����9@������@                      �?      �?      @      �?              �?                               @       @                      �?       @     pU@33333o}@                      �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff�7@     ��@      �?                              �?      �?              �?                                       @       @              �?       @fffffFV@fffffFV@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@      �?                              L@      �?       @      �?       @                       @       @       @              �?      @fffffVZ@3333s��@                      �?              3@      �?                                                                                      @33333sF@33333=�@      �?              �?             �I@      �?                       @       @       @       @       @       @       @      �?      �?fffff�T@����Ӱ@      �?              �?      �?      5@      �?       @      �?               @       @               @       @                       @�����Z@ffff�۠@      �?      �?                      B@      �?       @      �?       @                               @                      �?       @fffff�V@fffff�@                      �?      �?     �Q@      �?       @      �?       @       @       @               @               @      �?      �?     �X@ffff���@      �?                              L@      �?                       @               @                              �?              @�����YJ@fffff��@      �?                              G@      �?       @      �?               @       @       @       @       @       @               @�����)[@33333'�@      �?              �?      �?     @Q@      �?       @      �?               @       @               @              �?              �?     �W@    @o�@      �?              �?              �?      �?       @      �?                                                              �?        fffff�R@fffff�R@      �?      �?                       @      �?       @      �?                                                              �?      @fffff�R@����̌c@              �?                      @              �?                                               @       @                       @������F@     �h@      �?              �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�����9@33333��@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����L3@�����YK@                                     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�����:@������@                                      R@      �?       @      �?       @       @       @       @       @       @       @              �?33333�\@    �j�@      �?                              4@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @33333�3@fffff�y@      �?              �?             �I@      �?       @      �?               @                               @      �?      �?      �?fffff�V@���̌�@      �?              �?             @P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?ffffff4@������@      �?              �?              I@              �?               @                       @       @              �?      �?        �����9F@ffff��@              �?      �?              R@      �?       @      �?       @       @       @               @       @       @      �?       @�����\@�����n�@      �?      �?      �?      �?      R@      �?              �?       @               @       @       @       @       @      �?      �?fffffZ@3333��@                                     �B@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@fffffj�@              �?                      @      �?       @      �?                                                              �?      �?33333�R@     p@                                      =@      �?       @               @                                       @              �?       @fffff�P@�������@      �?      �?                       @      �?       @      �?                       @                                      �?       @     PT@�����O�@      �?      �?                      @@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@�����]�@      �?              �?      �?      7@      �?       @                       @               @                       @              @������M@������@      �?              �?      �?      R@      �?       @      �?       @               @               @       @      �?      �?        fffff�Z@    ���@      �?              �?      �?      Q@      �?              �?       @       @       @               @       @       @      �?             PZ@ffff&�@      �?                             �A@      �?       @               @               @                                      �?       @������M@�����]�@      �?      �?      �?             �@@      �?              �?       @       @               @               @      �?      �?       @33333cW@     ߧ@      �?      �?      �?      �?      =@      �?       @      �?                       @               @       @              �?       @������Y@�����)�@      �?              �?      �?      $@              �?               @       @       @       @               @       @              �?������J@     H�@                      �?              1@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����Y3@     0s@      �?      �?      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      @     �\@�����E�@      �?                              9@      �?       @               @       @       @       @               @                             pT@33333��@      �?              �?      �?      J@      �?                       @       @       @               @       @       @               @������S@�����`�@                                      @      �?              �?                                       @                      �?       @������S@����̔n@      �?                              $@      �?                                                                              �?      �?�����lF@fffff6{@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@     �3@                      �?             �M@      �?       @                       @               @       @       @      �?      �?       @fffffT@33333U�@      �?                              &@      �?                               @                       @              �?      �?       @     �N@�����φ@      �?                              ,@              �?                               @               @       @              �?       @     `I@     F�@                      �?      �?       @      �?              �?               @                       @                      �?       @33333�T@fffff@�@                      �?              4@      �?               @      �?      �?      �?      �?      �?      �?                             @3@     tw@      �?                              R@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?������3@     �@      �?                              *@      �?       @      �?                               @       @       @                       @     0Y@     ��@      �?                              �?      �?                                               @                              �?       @fffff�H@fffff�H@      �?      �?      �?              R@      �?       @      �?               @       @               @       @       @      �?        �����	Z@3333�	�@                      �?      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?       @                     �3@fffff>�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@33333�Z@              �?                       @              �?                               @                                      �?       @ffffff>@������S@                                      *@      �?               @      �?      �?      �?      �?      �?      �?      �?              @3333334@     q@      �?      �?      �?              O@      �?       @      �?               @                               @              �?        33333sV@���̌��@      �?      �?      �?      �?      &@      �?       @      �?                                                              �?      �?������R@fffff:�@      �?      �?                      .@      �?              �?               @                                              �?       @������R@33333ɐ@      �?              �?      �?     �Q@      �?       @      �?               @                       @       @       @                33333�X@    �˺@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y3@�����,G@      �?                              .@      �?       @                       @               @                              �?      �?�����LM@�����]�@      �?      �?      �?              C@              �?                                                                      �?       @������8@     ލ@      �?                              6@      �?       @      �?               @                       @       @              �?       @�����)Y@ffff�ߢ@              �?      �?      �?      �?      �?              �?                                                              �?       @     PQ@     PQ@      �?              �?      �?     �O@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     @9@33333��@      �?      �?                      (@              �?                               @       @               @              �?       @33333�E@�����w�@                                      B@      �?       @               @               @       @       @       @      �?      �?      �?�����iV@33333(�@      �?                              K@      �?       @      �?                       @                       @                      �?�����YV@    ��@      �?      �?      �?      �?     �N@      �?       @      �?               @                       @       @      �?               @     �X@����LQ�@                      �?              >@      �?       @      �?                                               @              �?       @     @U@    ���@              �?                      @      �?              �?                       @               @                      �?       @fffffU@33333�@                                      @      �?       @                                               @                      �?       @      N@     Pe@                                      �?      �?       @      �?                                       @       @              �?       @fffff�W@fffff�W@                                     �Q@      �?       @      �?               @       @       @                      �?      �?             �V@3333��@                      �?             �L@      �?       @                       @       @       @       @              �?                fffff�R@3333��@                                      E@      �?       @                               @       @       @       @       @      �?      �?����̜S@�����Z�@                                      1@      �?       @      �?       @       @                       @                      �?       @������W@     F�@                      �?      �?      H@      �?                       @       @       @                       @       @      �?      �?fffff�Q@�����L�@      �?              �?              R@      �?       @               @       @       @       @       @       @       @      �?        fffff�U@����V�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@                      �?              P@      �?       @               @       @       @       @               @       @      �?      @33333ST@����L	�@      �?                              ,@              �?                               @       @       @       @              �?       @     �K@������@      �?              �?      �?      3@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@33333[v@      �?                      �?      9@      �?              �?               @                       @       @              �?       @������W@    �!�@      �?                              (@      �?              �?                                       @                      �?       @�����\T@     ��@      �?                              (@      �?                       @                       @                                      @33333SL@�����v�@      �?      �?      �?              J@      �?              �?       @               @       @       @       @      �?      �?        �����Z@    @i�@      �?                               @      �?                                                                                      @33333SF@������R@                                      4@      �?               @      �?      �?      �?      �?      �?      �?              �?             �3@     �y@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @fffff&4@fffffvd@      �?                              @      �?       @      �?       @                                                      �?       @fffffT@fffffu@                                      @              �?                                               @       @                      �?     �F@33333�r@      �?                               @      �?       @      �?                                               @              �?       @33333�U@33333M�@      �?                              .@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@�����	s@      �?                               @              �?               @                                                      �?       @33333s>@fffffNl@                      �?              :@              �?               @               @                              �?              �?33333�A@����̔�@                                      H@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?      8@33333|�@                                     �J@      �?       @      �?               @       @               @       @       @               @33333cZ@    @2�@                                      "@      �?                               @               @       @                              @     �P@fffffd�@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @              �?�����,V@����Ye�@                      �?      �?      P@      �?               @      �?      �?      �?      �?      �?      �?       @              @3333334@     ��@      �?              �?              P@      �?       @      �?               @               @       @       @       @      �?       @     PZ@fffff��@                              �?       @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@33333sd@      �?              �?              $@      �?              �?                                       @                      �?       @������S@�����Ɋ@      �?              �?      �?      R@      �?       @      �?       @       @       @               @       @       @      �?      �?�����[@    @W�@              �?                      @              �?                                               @       @              �?       @333333F@�����pp@      �?              �?              8@      �?       @      �?                                       @       @              �?       @     @W@������@      �?                              $@      �?                       @                                                      �?      @33333�I@     d�@                                       @      �?                               @                       @                      �?       @     �M@������\@      �?                      �?      *@      �?                                                       @       @                      �?������P@     ��@      �?      �?      �?              B@      �?       @      �?                                               @              �?       @fffffU@33333��@      �?                              4@      �?       @      �?                       @               @                      �?       @�����,V@����̅�@                                       @      �?              �?                                       @                      �?       @�����)T@�����b@      �?                               @      �?                               @                                              �?      @fffff&I@     0W@                                      E@      �?                       @       @               @               @      �?      �?      @������P@    ���@      �?                              $@      �?                                                                                      @      G@������~@      �?              �?      �?      A@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?������3@fffff6�@                      �?              O@      �?                       @               @       @       @       @       @              @     @T@ffff�y�@      �?      �?                      ,@      �?       @      �?                                       @       @              �?       @fffff�W@33333�@      �?                               @      �?       @      �?               @                       @       @                       @fffff6Y@fffff��@      �?                              9@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �����L9@�����"�@                                     �G@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     @4@33333�@      �?      �?      �?              7@      �?       @      �?               @       @               @       @              �?       @�����Z@3333��@                      �?      �?      @      �?              �?                                               @                       @fffff6T@     �r@      �?      �?      �?              ;@      �?       @                       @       @       @       @       @              �?        333333U@�����@      �?                             �L@      �?                       @               @               @       @       @      �?        fffff�R@����Yݰ@                                      =@      �?       @                       @                                      �?      �?       @     �K@�����P�@                                      *@      �?                       @                               @       @              �?       @������Q@�����ތ@                                      1@      �?               @      �?      �?      �?      �?      �?      �?       @              @ffffff3@�����`v@                      �?      �?      0@      �?              �?               @                                                             PR@     ��@                                      &@      �?                                       @       @                      �?                fffff�J@fffff\�@              �?      �?      �?     @P@      �?       @      �?               @       @               @       @      �?      �?       @������Z@    ���@                                      E@              �?               @       @       @       @               @      �?      �?       @     `K@ffff�X�@                                     �A@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����L7@������@                                      ,@      �?                                               @       @       @              �?       @�����iQ@33333ˌ@      �?                              =@      �?       @                       @       @                       @      �?              �?������Q@fffff��@                      �?              H@      �?       @      �?               @               @       @       @              �?      �?fffffFZ@���̌۳@      �?      �?      �?             �B@      �?       @      �?                                       @                      �?       @�����lU@����Lƨ@      �?                             �P@      �?              �?               @       @               @       @                       @     �X@    �6�@      �?              �?      �?      $@      �?       @       @      �?      �?      �?      �?      �?      �?              �?      @ffffff8@����̼o@              �?      �?              Q@      �?       @      �?               @                               @              �?        ffffffV@������@      �?                             �M@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        3333334@33333��@                      �?      �?      $@      �?               @      �?      �?      �?      �?      �?      �?              �?        ������3@     �h@              �?                       @      �?              �?                       @               @       @              �?      �?����̜W@�����7�@      �?              �?             �Q@      �?                       @               @       @       @       @       @      �?       @33333�T@ffff�ȶ@      �?                              @      �?       @      �?                                       @       @                      @     �W@     |�@      �?              �?      �?      O@      �?       @      �?       @       @                       @       @              �?       @     `Z@33333W�@      �?                              9@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?fffff�3@������@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@������[@                      �?              Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?33333�8@�����;�@                                      "@      �?       @      �?                                                              �?       @fffff6S@fffff��@      �?              �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������9@�����@�@      �?                             �B@      �?       @      �?               @               @       @       @      �?      �?      �?      Z@     ��@                      �?             �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @ffffff8@�����'�@      �?              �?      �?      6@      �?              �?               @       @               @       @      �?      �?      @33333Y@    �T�@      �?      �?      �?             �Q@              �?                       @       @               @       @              �?        fffff&J@����j�@                                     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ������9@fffff��@              �?                      0@      �?              �?                               @       @       @              �?       @����̜W@����̜�@                                       @      �?       @      �?                                                              �?       @     `R@�������@                      �?      �?     @Q@      �?       @      �?               @               @               @       @      �?        33333SW@������@                                       @      �?       @      �?                                                                      �?������R@�����db@                      �?      �?      R@      �?       @               @       @       @       @                       @      �?        ����̜Q@3333�-�@      �?                              4@      �?                       @               @                       @                      �?�����P@fffffڕ@                      �?             �Q@      �?       @                       @       @       @       @       @       @      �?        333333U@���̌�@                              �?      3@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@������x@                                       @      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�4@333333a@      �?                              Q@      �?       @      �?       @       @       @               @              �?                fffffVY@    �ƻ@      �?      �?                      �?      �?                                                                                       @      F@      F@                      �?      �?     �H@      �?       @      �?               @                       @       @              �?       @fffff�X@33333�@      �?              �?              =@      �?       @      �?       @       @                                              �?       @�����U@33333F�@                                      ?@      �?              �?       @               @       @                                       @fffff�U@    �H�@      �?                              @      �?       @      �?                                                                       @ffffffR@     @�@      �?              �?      �?      Q@      �?       @      �?       @       @       @               @       @       @      �?       @����̌[@    �+�@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@������R@                      �?      �?      >@      �?                       @                       @               @                        33333�P@     �@                                      H@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                �����Y8@����̶�@      �?              �?             �G@      �?       @      �?                                       @       @      �?      �?      �?������W@     ӱ@                      �?      �?      8@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @33333�8@     ށ@              �?                     �D@      �?       @      �?               @       @               @       @              �?       @�����Z@3333�%�@      �?              �?              M@              �?                                               @       @      �?      �?      �?     �F@3333��@                      �?              J@      �?       @      �?               @       @               @       @              �?       @33333CZ@�������@      �?      �?                      8@      �?       @      �?               @       @               @       @              �?      �?����̼Y@fffff��@              �?                      F@      �?                                       @       @       @       @      �?                fffff�R@������@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @3333334@3333334@                                      @      �?              �?               @                                              �?        �����)S@������t@      �?              �?              8@      �?                       @                       @                                      @������J@fffff��@      �?                              $@      �?       @      �?                                                                       @33333�R@fffff��@      �?              �?              L@      �?       @      �?               @               @       @       @      �?      �?       @     �Z@����L��@      �?                              $@      �?       @      �?               @                                              �?        �����,T@fffff��@                              �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@333333X@      �?      �?                      @      �?              �?                                       @                      �?       @������S@�����@                      �?      �?      2@      �?               @      �?      �?      �?      �?      �?      �?              �?      @     @4@33333y@                                      �?              �?                                                                              @ffffff8@ffffff8@                                      $@      �?                                                                                      @     �F@33333�z@      �?              �?      �?      *@      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@     �o@                              �?      @      �?              �?                                                              �?       @33333�Q@fffff�}@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?              :@�����[�@      �?              �?      �?     �Q@      �?       @               @       @       @       @       @       @       @      �?      �?������V@����]�@      �?              �?              <@      �?       @      �?               @       @               @                              �?fffff&X@3333���@      �?      �?                      @      �?              �?                                                              �?       @������Q@�����]r@      �?              �?              6@      �?                       @                       @                              �?       @�����K@������@      �?      �?      �?              7@      �?       @      �?                                               @                       @33333�U@fffffߞ@      �?                      �?      "@      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@33333g@      �?              �?      �?     �M@      �?                               @       @       @       @       @      �?              �?     0S@ffff潱@              �?                     �F@      �?       @      �?                       @               @       @      �?      �?        ������Y@����Y�@                              �?      H@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@�����E�@                                      L@      �?       @      �?               @               @       @       @              �?        �����\Z@3333��@                                      @      �?       @      �?       @                                                      �?      @������S@������@      �?      �?      �?              8@      �?       @      �?               @       @               @       @              �?       @     Z@������@                                      $@      �?              �?                                               @              �?             T@     p�@                      �?              P@      �?              �?       @                       @       @       @      �?      �?      @�����9X@����Y��@                      �?      �?     �@@      �?       @      �?       @               @               @       @      �?      �?      @������Y@     �@                      �?              2@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@     (w@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                      9@     d�@                      �?      �?      ,@      �?       @      �?                                       @                      �?       @333333U@�����ϒ@                      �?      �?      N@              �?                       @                       @       @              �?       @     �H@ffff���@                      �?             �Q@              �?                               @       @               @       @      �?       @fffff�G@33333�@                      �?              :@      �?                               @       @               @       @       @      �?      �?     `R@�����Ɲ@      �?              �?      �?      2@      �?               @      �?      �?      �?      �?      �?      �?      �?                �����4@fffff�u@                      �?              F@      �?       @      �?                                       @       @              �?       @fffffX@�����@      �?                              8@      �?                       @       @               @                                        �����9N@     ��@                                      (@      �?               @      �?      �?      �?      �?      �?      �?                      @�����L4@fffff�n@                                      0@      �?               @      �?      �?      �?      �?      �?      �?      �?                �����4@������s@      �?              �?      �?      F@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?             �4@fffff�@                      �?              :@      �?               @      �?      �?      �?      �?      �?      �?      �?              @3333333@������|@                                      9@      �?                       @                       @       @       @              �?      �?�����	S@�����#�@                      �?              "@      �?              �?                                               @              �?       @     �S@������@                                      2@      �?                                       @                                      �?      @      I@������@                      �?             �K@      �?       @      �?               @                                              �?      �?     pS@fffff��@      �?                              =@      �?       @      �?                                               @              �?       @�����9U@fffff��@      �?              �?      �?      @      �?                               @       @                                      �?      @33333L@�����e@                                      $@      �?       @      �?               @                                              �?      �?     @T@fffff��@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�4@fffff�c@      �?                             �C@      �?              �?       @               @               @       @       @      �?       @�����Y@fffff��@                      �?      �?      7@      �?                       @       @               @                      �?      �?      @     �L@fffff�@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     �8@�������@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @������4@33333SN@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������3@33333}�@                      �?              6@      �?       @               @                       @       @       @              �?       @������S@     ;�@                      �?      �?     �Q@      �?                       @               @               @       @       @              �?33333cS@����YƵ@                                      @      �?              �?                                       @       @              �?       @�����\V@fffffn@              �?                      L@      �?       @      �?               @       @       @       @       @      �?      �?       @������[@ffff��@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?     @8@������@                                     �L@      �?       @      �?       @       @               @                              �?        33333�U@������@                                      0@      �?              �?               @                               @              �?       @     �U@fffff�@      �?                              $@              �?                       @               @                                       @     �A@�����\x@      �?                              :@      �?       @      �?       @       @                                              �?      �?������U@    �A�@              �?      �?               @      �?                               @                                                      �?33333I@fffff�\@              �?                      @      �?              �?                                       @                      �?       @fffff�S@�����Lr@              �?      �?              N@              �?                       @                       @       @       @      �?      �?������H@������@      �?              �?      �?      E@      �?                       @                       @               @      �?              �?������O@3333���@      �?              �?      �?     �@@      �?                                       @       @       @       @      �?      �?      @�����yR@����ʢ@                      �?      �?     �C@      �?              �?                       @       @                              �?             `T@�����F�@      �?                      �?      @      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @ffffff:@     P^@                                      �?      �?              �?                                       @                               @33333�S@33333�S@      �?                              2@      �?       @      �?                                                              �?        fffff�R@33333̕@      �?                              �?      �?              �?                                                              �?       @33333�Q@33333�Q@                                      "@              �?               @               @       @       @       @                      @     @M@�����ހ@      �?              �?      �?      R@      �?       @      �?       @       @       @               @       @       @      �?        33333�[@ffff��@      �?              �?               @      �?                               @       @                                      �?      @     `K@������{@              �?                      E@      �?       @      �?               @       @               @       @              �?             0Z@3333s�@      �?              �?      �?     �Q@      �?       @      �?       @                               @       @       @      �?       @�����LX@����L��@      �?                              :@              �?                               @       @                                       @     �A@     �@      �?                              �?      �?       @                                                                      �?      �?fffff�H@fffff�H@      �?              �?              B@      �?               @      �?      �?      �?      �?      �?      �?      �?                ������4@fffff��@      �?                              :@      �?                                                                                       @������F@�����D�@      �?              �?              H@      �?               @      �?      �?      �?      �?      �?      �?       @              @     @3@����̸�@                      �?             �F@      �?       @      �?       @       @       @       @       @       @      �?              @33333S\@    @��@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@33333s]@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@     �O@                                       @      �?               @      �?      �?      �?      �?      �?      �?              �?      @����̌4@������@@      �?                               @      �?                                                                              �?       @33333�F@     �X@      �?                              @      �?       @      �?               @       @               @       @              �?        fffffVZ@     4t@                                      B@              �?               @       @       @       @               @       @      �?      @����̌J@     ��@      �?              �?              D@      �?       @      �?                                       @       @              �?        fffffFX@ffff���@                                      @      �?              �?                                               @              �?       @33333�S@33333Y�@                                     �C@      �?              �?                       @       @                       @      �?       @�����T@�����@      �?                              :@      �?       @      �?                       @       @                              �?      @33333U@33333ӡ@      �?              �?      �?     �C@      �?                       @               @       @       @       @      �?              �?      T@ffff�ݨ@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@                                      >@      �?              �?                               @       @                               @�����IU@�������@      �?              �?      �?      @      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�����8@fffffFR@                                      ;@      �?               @      �?      �?      �?      �?      �?      �?       @      �?             @4@�����р@              �?                      .@      �?       @                                       @                                      �?     �K@����̨�@                      �?      �?       @      �?                       @       @                                                      @33333SK@     $~@      �?      �?      �?      �?     �D@      �?       @      �?               @       @       @       @       @      �?      �?       @������[@ffff涱@      �?                              ;@      �?       @                               @       @                                       @������M@�����.�@      �?              �?              J@      �?              �?       @       @       @       @       @       @       @      �?       @33333�Z@     o�@      �?              �?      �?     �J@      �?       @               @       @                               @       @                �����lQ@����̬@      �?      �?                      "@      �?              �?                                               @              �?       @33333�S@ffffft�@      �?                              0@      �?       @                       @       @                       @              �?        ������Q@fffff�@      �?              �?      �?     �O@      �?       @               @               @       @               @       @              @������R@3333�D�@      �?                              @      �?              �?                                               @              �?       @fffffT@������o@                              �?      8@      �?               @      �?      �?      �?      �?      �?      �?      �?                �����5@fffff��@      �?              �?      �?      0@      �?       @               @       @               @       @       @                       @�����9U@     ٕ@                                      @      �?              �?                       @                       @                       @������T@�����@      �?                              3@              �?                               @               @                      �?       @33333�C@������@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�3@fffff�3@      �?              �?              4@      �?                       @                       @               @      �?      �?      @�����	P@������@                      �?      �?     �@@      �?       @      �?                                               @                      �?������U@fffffs�@              �?      �?              M@      �?              �?       @       @               @       @       @      �?      �?      �?     `Z@    �=�@                                      @              �?                               @               @       @              �?       @������G@�����s@                                      H@      �?                       @               @       @                      �?      �?      �?�����,N@����̠�@      �?              �?      �?     �M@      �?                       @       @       @       @       @       @       @      �?       @     �U@     B�@                                      "@      �?       @      �?                                       @       @              �?       @     �W@33333ϋ@      �?                              J@      �?       @      �?                       @                       @       @      �?      �?�����\V@    ��@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?       @              @33333s4@33333s4@              �?                      P@              �?                       @               @       @                      �?       @������E@     ~�@                                     �H@      �?                                       @       @       @       @       @      �?        ����̜R@������@      �?                             �A@      �?       @      �?                                                                      �?fffff�R@������@                                      3@      �?                                                               @              �?       @�����L@������@      �?      �?                      (@      �?       @      �?                                                              �?      �?33333SR@fffff��@      �?              �?      �?      ;@      �?       @      �?                                                              �?             �R@     $�@                      �?      �?     @Q@      �?       @               @               @       @                       @      �?      �?�����	P@������@                      �?              @@      �?              �?       @                                                      �?             �R@fffff)�@      �?                      �?      N@      �?       @               @               @       @       @       @       @      �?       @�����<U@�����x�@                      �?      �?      F@      �?                       @                       @                                              L@�����@      �?                              5@      �?       @      �?                                                                      @33333�R@����̊�@              �?      �?              =@      �?       @      �?                       @               @       @              �?        33333�X@3333��@      �?              �?             �K@              �?                               @       @       @       @              �?        fffffFK@�����D�@      �?                              (@      �?       @      �?                               @       @       @              �?      @������X@     ��@                                      @              �?                                                                      �?      @     @8@33333X@                                      �?              �?                                       @                                      @����̌>@����̌>@                      �?              @      �?       @      �?               @                               @              �?       @     �V@     �@                      �?             �Q@              �?                       @       @       @       @       @       @      �?      �?33333�N@����Yְ@                      �?              P@      �?       @                               @       @                      �?                �����,M@ffff�X�@                      �?      �?     �N@      �?       @               @       @                                                       @fffff�M@     s�@                                       @      �?              �?               @                       @                      �?        ������U@     �f@                                      @      �?               @      �?      �?      �?      �?      �?      �?                       @����̌3@fffff�N@                      �?              G@      �?                               @               @       @               @      �?      �?�����P@     ��@                                      A@      �?                       @               @       @       @       @      �?      �?        ������S@�����N�@              �?                      @              �?                       @                                                       @33333s<@�����a`@      �?              �?              R@      �?       @               @       @       @       @       @       @       @              �?33333W@ffff�?�@      �?              �?      �?      @              �?               @       @       @                               @              @fffffFC@     �q@      �?              �?              @      �?               @      �?      �?      �?      �?      �?      �?                              4@33333�H@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                       @����̌4@����̌4@              �?                      @      �?              �?                       @               @                      �?      @fffff6U@������y@                                      3@              �?                       @                               @              �?       @������C@fffff0�@      �?      �?                      �?              �?                       @       @                       @              �?       @fffff�E@fffff�E@                      �?      �?      @@      �?                       @       @               @                                        33333�N@�����"�@      �?      �?                      4@      �?              �?                                                                      �?33333�Q@����̴�@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?33333s:@     �@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����8@�������@      �?                              "@      �?              �?                                               @              �?       @333333T@�����H�@      �?                              (@      �?       @      �?                                       @                      �?       @�����U@33333��@      �?                              @      �?              �?                                       @                      �?       @fffff&T@������y@                                      @      �?              �?                                                                      �?33333�Q@33333{@      �?              �?             �L@      �?       @      �?                       @       @       @       @       @               @������Z@�����Q�@                      �?      �?      P@      �?       @      �?       @       @               @       @       @       @                33333�[@����LU�@      �?                             @Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����L3@�������@                                      @              �?                                               @                              �?������A@�����<[@      �?              �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @                3333334@     ��@      �?              �?      �?      :@      �?              �?                                               @      �?                ����̼S@     ɟ@                                      &@      �?                                       @       @               @      �?              �?�����9P@     ʅ@      �?              �?      �?      0@      �?               @      �?      �?      �?      �?      �?      �?                       @     �3@fffff�s@              �?      �?      �?      O@      �?       @      �?               @       @                       @              �?      �?fffffX@����Y��@              �?                      �?      �?              �?                                                              �?       @     �Q@     �Q@      �?                              $@      �?               @      �?      �?      �?      �?      �?      �?                      �?      4@fffff�h@      �?                              "@      �?              �?                       @               @       @              �?       @33333�W@33333]�@                      �?             �P@      �?       @      �?       @       @               @                      �?               @     @V@�����
�@                                      9@      �?       @               @       @       @       @       @                      �?        fffff�S@�������@      �?                              2@      �?       @               @                                                              @      L@�����N�@                      �?      �?      ;@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����̌4@fffff:�@      �?      �?                      C@      �?       @      �?                                       @       @                       @     �W@     ��@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @3333333@3333333@                                      (@      �?              �?                                               @                        fffff�S@fffff��@                                     �Q@      �?       @               @       @       @               @       @       @              @�����,U@����g�@      �?                      �?      �?      �?              �?                                                                             pQ@     pQ@                                      9@              �?                               @               @       @              �?       @      H@333337�@                              �?      �?      �?              �?                                       @       @              �?       @fffffVV@fffffVV@              �?                      5@      �?       @      �?                                       @       @              �?       @     �W@     מ@                                      �?      �?              �?                                                              �?       @fffff�Q@fffff�Q@                                      &@      �?       @      �?                               @       @                               @������V@�����ߎ@      �?      �?                      3@      �?              �?       @                                       @              �?       @33333�U@33333��@      �?              �?              @@      �?       @               @                       @       @              �?      �?      �?333333R@����:�@                              �?      @      �?       @      �?               @       @                                                33333U@������t@                      �?             �@@      �?              �?       @               @       @       @       @      �?      �?       @     �Y@����B�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?     �4@fffff�P@                                      7@      �?       @      �?                                       @       @              �?       @     `W@����K�@                      �?              @      �?              �?                                                              �?        �����LQ@������}@      �?      �?                       @      �?       @      �?                                                              �?      @fffff&R@�����Ic@      �?              �?      �?      Q@      �?              �?               @       @       @       @       @      �?              �?     pZ@    ���@      �?              �?      �?      �?      �?              �?                                               @                       @      T@      T@      �?      �?      �?              R@      �?       @                       @       @       @       @               @              �?fffffVS@    @�@                      �?              @      �?       @                                                                               @�����,I@����̨s@      �?                      �?      F@      �?               @      �?      �?      �?      �?      �?      �?       @                ����̌3@�������@              �?                      �?      �?              �?                                       @       @              �?       @33333SV@33333SV@      �?                      �?     �E@              �?               @       @       @                                      �?       @�����9D@fffff�@                      �?      �?      E@      �?       @       @      �?      �?      �?      �?      �?      �?       @               @33333�6@     ��@      �?      �?      �?              R@              �?               @       @       @       @       @       @       @      �?      �?�����P@����!�@      �?                             @P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �9@     ۙ@      �?              �?              =@      �?              �?                       @                                      �?      �?33333�R@����̮�@                                      �?      �?              �?                       @                                                     `R@     `R@      �?              �?              2@      �?       @                       @                                                      �?ffffffL@�����ʐ@      �?              �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����4@     A�@                                      "@      �?              �?       @                                                      �?       @fffff�R@�����!�@      �?              �?             �G@      �?       @      �?               @       @                                      �?        fffff�T@     ¯@                      �?      �?      �?      �?              �?                                                              �?      @fffffFQ@fffffFQ@      �?              �?      �?      9@      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff&3@������}@                                      $@      �?       @      �?                               @       @       @              �?       @     �X@     ��@              �?                      D@      �?              �?                                       @       @              �?       @33333�V@33333��@                      �?              N@              �?               @       @               @                       @                ������B@fffff�@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?       @     �\@ffff&��@                      �?              C@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?     @4@     v�@                              �?       @      �?       @      �?       @                                                              �?33333#T@33333�g@                                      (@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����L3@     �l@      �?                              >@      �?       @      �?       @       @       @       @                              �?      �?     �W@�����H�@      �?              �?      �?      L@      �?       @       @      �?      �?      �?      �?      �?      �?       @                fffff&8@     �@                      �?             �P@      �?       @      �?       @               @       @       @       @      �?      �?       @     �[@ffff�W�@                      �?             �Q@      �?       @      �?       @               @               @       @      �?      �?      �?fffffZ@    @��@                      �?      �?      >@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�����9@fffff��@      �?      �?      �?              R@      �?       @      �?               @       @       @       @       @       @      �?        ������[@�����V�@                      �?      �?      (@      �?       @      �?               @       @                                      �?       @      U@33333��@                                      (@              �?               @                       @                      �?      �?      @������@@333337{@                      �?      �?     �M@      �?               @      �?      �?      �?      �?      �?      �?       @              @������4@     �@                      �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @                �����4@fffffӖ@                      �?      �?     �H@              �?               @                       @                      �?      �?      �?fffff�A@     ؛@                      �?      �?      @      �?                                                       @                               @�����lK@�����1v@              �?                       @      �?       @      �?                               @       @       @              �?      �?�����	Y@fffffd�@      �?              �?             �K@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333�9@�������@      �?                             �G@      �?       @      �?               @       @               @       @      �?      �?       @fffff�Y@����L�@      �?                             �E@      �?       @      �?               @                                              �?       @fffffvS@3333�K�@      �?      �?      �?              �?      �?       @      �?                                       @       @              �?       @fffff�W@fffff�W@      �?              �?      �?     �B@              �?               @               @       @                      �?      �?       @�����D@fffff՗@      �?              �?      �?      I@      �?       @      �?               @               @       @       @                       @������Y@����ϳ@      �?              �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@     ѕ@      �?                             @Q@      �?       @      �?               @       @       @       @               @      �?      �?�����iX@���̌W�@      �?                              @      �?       @                                                                              �?     �I@33333#i@      �?                              "@      �?       @      �?       @                                                      �?       @�����IT@�������@                      �?              9@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      @������:@fffff�@                                     �D@      �?              �?                                                                             �Q@����h�@      �?      �?      �?              0@      �?              �?               @                                              �?      �?33333�R@     i�@      �?                              M@      �?               @      �?      �?      �?      �?      �?      �?       @              @������4@     �@                                     �M@      �?              �?                       @               @       @       @               @33333�W@3333s�@                      �?              6@      �?              �?                                                              �?       @     PQ@     H�@      �?                              @      �?                       @               @               @       @              �?       @�����YS@������i@                                      (@      �?       @      �?                                               @              �?       @33333�U@�������@                                      ?@      �?       @      �?       @               @                                      �?      �?     0U@�����j�@                                     �D@      �?       @                               @       @               @      �?      �?       @fffff&Q@����z�@      �?              �?      �?      3@      �?       @      �?                       @       @       @       @                       @33333�Y@�����r�@                                      "@      �?                                               @       @                      �?             �M@fffff��@                                     �L@      �?       @      �?               @               @               @      �?               @����̬W@3333�\�@                      �?              @@      �?              �?               @                               @                        �����	U@ffff�3�@      �?      �?                      "@      �?       @      �?                                               @              �?      �?�����U@     �@                      �?      �?     �A@      �?       @               @       @                                              �?      �?������M@����̱�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      �?�����L3@�����L3@                      �?      �?     �P@      �?                       @       @               @                       @      �?      �?�����M@�����ŭ@      �?              �?      �?      G@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�����4@�����F�@      �?      �?      �?              $@      �?       @      �?                       @                       @              �?       @33333sV@fffff��@                                      ?@      �?       @      �?                               @                              �?      �?fffff�S@����LȢ@      �?                             �B@      �?       @      �?       @                               @                      �?       @������V@    �R�@                                     �O@      �?       @      �?               @       @       @       @       @              �?      �?fffffv[@3333�Z�@                      �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����Y4@33333�t@                                      $@              �?                                       @                       @      �?      @������=@����̰r@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                       @33333�3@33333�3@                                      @      �?       @      �?               @               @               @              �?       @     `W@33333�v@      �?                              6@              �?                               @       @       @       @       @                     `L@fffffc�@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@33333C@      �?                      �?       @              �?                                                                              @     �9@fffff�j@                      �?              G@      �?                       @       @               @               @      �?              @fffff�Q@����>�@      �?                              F@      �?       @      �?       @       @       @               @       @              �?       @     �[@ffff&3�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����4@                                      $@      �?       @      �?                                               @                       @����̜U@�������@      �?              �?      �?      =@              �?               @       @       @       @               @      �?      �?      �?����̬K@����̓�@                      �?      �?     �A@      �?       @               @               @       @       @                               @     R@�����@              �?                      0@      �?       @      �?                                       @       @              �?       @�����	X@������@                                       @      �?                                       @       @       @       @                       @�����S@�����d@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@33333�d@      �?              �?              >@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����3@fffff�@                              �?       @      �?       @      �?                                       @       @              �?        ����̌W@�����9h@      �?                              �?      �?                       @                                                              @     �I@     �I@                      �?      �?     �B@      �?       @       @      �?      �?      �?      �?      �?      �?                      @33333s:@�����|�@                                      C@      �?       @               @       @       @               @       @      �?                fffffU@����L�@      �?              �?      �?      2@              �?                       @       @               @              �?              �?333333G@33333c�@      �?              �?              4@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�4@     z@      �?                              3@      �?       @                               @       @                                       @fffff�M@fffff�@      �?                             �H@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?fffff�3@������@      �?      �?      �?      �?     �A@      �?                               @               @       @       @              �?       @33333S@fffffv�@                                       @      �?       @      �?       @                       @       @       @              �?        fffff�Y@fffffz�@                      �?      �?      R@      �?                       @       @       @               @               @      �?      �?������Q@ffff&��@      �?              �?      �?     �Q@      �?       @      �?               @                       @       @      �?                33333#Y@    �ɻ@      �?                              0@      �?       @                       @                                                       @fffff�K@�����Z�@                      �?      �?      6@      �?               @      �?      �?      �?      �?      �?      �?                        �����3@�����`|@                      �?      �?       @      �?              �?                                                                       @������Q@�����db@              �?      �?             @P@      �?       @      �?               @       @               @       @              �?        333333[@3333s��@      �?              �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����Y9@33333ޜ@      �?                              �?      �?                                                       @       @              �?      @ffffffO@ffffffO@                      �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����L4@�����j�@                              �?      �?      �?              �?                                       @                      �?       @fffff�S@fffff�S@      �?      �?      �?              4@      �?       @      �?                                       @       @              �?       @33333�W@�������@                                      �?      �?              �?                                                                       @fffff�Q@fffff�Q@      �?                              4@      �?       @      �?                                       @                      �?       @     PU@     �@      �?      �?      �?              O@      �?       @      �?       @       @       @                                      �?       @fffffFV@����L�@      �?                              @      �?       @      �?                                               @              �?      @�����LU@fffffԂ@      �?              �?             �H@      �?              �?                       @       @       @       @      �?      �?      �?     �X@�����8�@      �?                      �?     �G@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?����̌4@fffff��@                      �?      �?     �L@      �?                       @                               @       @      �?      �?        fffff�Q@�������@                                      �?      �?                       @       @                                              �?       @33333sK@33333sK@      �?                             �O@      �?       @               @       @       @       @                      �?                333333Q@����Y�@                      �?      �?     @P@      �?       @      �?       @               @               @       @       @      �?      �?33333Z@����LE�@              �?                      &@      �?       @      �?                                               @              �?      �?333333U@�����V�@                      �?      �?     �N@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����3@33333ߑ@      �?                              �?      �?                       @                                                      �?      @fffffFH@fffffFH@      �?                              �?      �?              �?       @                                       @              �?      @fffff&U@fffff&U@      �?              �?              5@      �?       @      �?               @       @       @       @       @              �?       @������[@33333�@                                      @      �?              �?                               @               @                       @33333sU@33333q@      �?      �?      �?              @      �?       @      �?                       @                                      �?        ������S@33333u@      �?      �?      �?      �?      �?      �?                                               @                              �?      �?     �H@     �H@                                      5@      �?              �?               @               @       @       @              �?        ������X@�������@      �?                              .@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @�����Y:@������w@      �?                              �?      �?       @                       @                                                       @fffff&K@fffff&K@                      �?              L@      �?       @      �?               @                       @       @      �?      �?       @     �X@����Y��@      �?              �?              @      �?       @      �?       @                                       @              �?       @�����IV@     �y@                                      �?      �?                                                                                      @������F@������F@      �?                              @              �?                       @               @                              �?      @�����lB@�����,[@      �?              �?              �?      �?              �?                                                                       @     �Q@     �Q@              �?      �?              @      �?              �?                                                              �?       @fffffVQ@�����Yu@                      �?      �?      ,@      �?              �?                                               @              �?        �����9T@33333�@      �?              �?      �?      E@              �?               @               @       @       @               @              �?33333H@33333��@                                     �C@      �?              �?       @               @       @       @              �?      �?       @33333�W@3333�٬@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@     �3@                                      7@      �?                                       @                                              �?������H@     �@                                      N@      �?               @      �?      �?      �?      �?      �?      �?       @                ������3@fffff��@      �?                      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������3@33333J�@                                     �I@              �?                       @       @               @       @      �?      �?      �?333333L@     �@      �?      �?              �?      �?      �?                                       @                                      �?      @33333I@33333I@                                      4@      �?              �?       @               @               @                      �?        �����YV@�����<�@                      �?              N@      �?       @      �?               @       @               @       @              �?       @������Z@    @�@                                      M@      �?       @               @       @       @       @                      �?      �?      �?fffff�Q@33333˰@      �?      �?      �?              G@      �?       @      �?                       @               @       @              �?       @fffff�X@ffff�Ա@                      �?              R@      �?       @      �?               @                       @       @       @      �?      �?�����lX@3333�պ@      �?              �?              R@      �?       @      �?       @       @       @                       @       @      �?       @������X@������@                      �?              *@      �?       @      �?               @       @               @                               @fffff�W@fffff��@                                      �?      �?                                                       @                      �?      �?     �K@     �K@      �?                              @      �?                               @               @               @              �?        ffffffP@fffff>u@      �?      �?      �?             �I@      �?       @      �?       @               @               @                      �?        33333sW@3333�@                                      ;@      �?                               @       @       @       @       @      �?              @����̌S@ffff�=�@      �?              �?      �?      7@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�4@     `|@                      �?              &@      �?                                                                              �?       @fffffF@33333;~@      �?                               @      �?                                               @       @       @                       @33333�Q@����̌`@                                      (@      �?                                                                                        fffff�E@������@                                      1@      �?       @       @      �?      �?      �?      �?      �?      �?                      @������8@     �}@      �?                              Q@      �?       @               @       @       @                       @      �?      �?      �?�����9S@     ��@      �?                              *@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @33333�3@������o@                      �?             �L@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ������3@     ��@      �?                              H@      �?                               @       @       @       @       @       @              �?������S@     w�@              �?      �?             �B@      �?       @      �?                                                              �?       @      S@����Lh�@                                      K@      �?       @      �?       @               @               @       @      �?      �?        ������Y@�����@      �?                      �?      4@      �?               @      �?      �?      �?      �?      �?      �?              �?       @ffffff3@     hw@              �?      �?              K@      �?       @      �?               @                       @       @      �?      �?      �?     `Y@������@      �?                              @      �?                                       @       @       @       @              �?       @������R@33333�r@                      �?      �?      R@              �?               @       @       @       @               @       @              �?33333�K@����P�@      �?                              &@      �?              �?       @                                                      �?       @     `R@     ��@                                      @      �?                       @       @               @       @       @              �?       @     �S@fffff؁@                      �?      �?     �B@      �?       @      �?                                       @       @              �?       @     �W@����L�@      �?              �?      �?      O@      �?               @      �?      �?      �?      �?      �?      �?      �?                33333�3@33333s�@              �?      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?     0]@ffff�*�@      �?                              ,@      �?       @      �?                               @       @                      �?       @�����|V@�����i�@      �?              �?      �?     �B@      �?               @      �?      �?      �?      �?      �?      �?       @                ������3@����̰�@      �?              �?      �?      >@      �?       @               @       @       @       @                                       @fffff�P@�����@�@                                      F@      �?       @      �?               @       @                                      �?        333333U@����-�@      �?                             �G@      �?                       @       @       @       @       @       @      �?      �?        ����̼U@ffff�*�@      �?                             �Q@              �?               @       @       @       @       @               @                ������J@����La�@      �?      �?                     �K@              �?                               @               @       @      �?      �?        fffffI@ffff�n�@              �?                     �G@      �?       @      �?               @               @       @                      �?       @33333�W@���̌��@      �?                              P@      �?              �?       @       @                       @       @      �?      �?      �?33333Y@�����˹@      �?              �?      �?      R@      �?                       @               @       @       @       @       @      �?       @333333T@���̌`�@      �?              �?      �?      �?      �?              �?                                                              �?      @������Q@������Q@                      �?               @      �?                                                                              �?       @     �F@     pV@                                     �P@              �?               @               @       @       @       @       @      �?        ����̬N@fffffa�@      �?              �?      �?      >@      �?       @      �?                                       @                               @�����\U@ffff曣@      �?                              �?      �?       @                                                                      �?       @33333I@33333I@      �?                               @      �?       @      �?                                               @              �?       @     �U@fffff�d@              �?                      B@      �?       @      �?                                                              �?        ������R@ffff�Ƥ@                      �?              7@      �?                       @               @       @               @      �?      �?             0Q@�����e�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @3333334@3333334@                                      @      �?              �?                       @                                      �?       @������R@     h�@      �?              �?              F@      �?                               @       @       @       @              �?      �?       @����̼Q@ffff�d�@                      �?      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @fffff�8@     A�@      �?                              3@      �?              �?               @                                              �?      �?fffffvR@     B�@      �?              �?      �?      J@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @������8@fffff4�@      �?                              @      �?                                               @                              �?       @������H@�����k@                                       @      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@     �C@      �?                              O@      �?       @      �?                       @               @       @      �?      �?       @     0X@fffff�@      �?                              M@      �?              �?       @       @                       @       @      �?                ������X@3333�X�@      �?                              �?      �?       @      �?                                                              �?       @33333�R@33333�R@      �?              �?      �?     @Q@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff�\@������@      �?                              �?      �?                                                                                      @333333F@333333F@      �?              �?      �?      ;@      �?       @      �?               @               @                              �?      �?�����LU@33333Ϡ@                                      N@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @      9@33333��@                      �?      �?      R@      �?       @               @               @       @                       @                fffff�P@����̖�@              �?      �?              H@      �?                               @                               @      �?      �?        �����yM@fffff˥@              �?      �?             �A@      �?       @      �?       @       @               @       @                      �?              Y@3333���@      �?              �?      �?      >@      �?       @      �?       @       @                       @                      �?       @������W@fffff-�@                      �?             �G@      �?       @      �?       @       @       @               @                      �?       @     �X@3333���@              �?      �?             �Q@      �?       @      �?               @               @       @       @       @      �?        �����Z@����Y��@      �?      �?                       @      �?              �?                                                              �?       @�����lQ@����̆�@      �?                              :@      �?                                               @                                        33333�H@33333U�@      �?                              K@      �?              �?       @       @               @       @       @      �?      �?      �?�����YZ@fffff�@              �?                     �D@      �?       @      �?       @       @       @               @       @              �?       @�����L\@    �Q�@                                      *@      �?       @               @               @               @       @              �?       @     �S@������@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @                ������3@�����֕@                      �?      �?      ?@      �?               @      �?      �?      �?      �?      �?      �?              �?      @����̌3@�������@      �?              �?      �?     �I@      �?               @      �?      �?      �?      �?      �?      �?       @              �?����̌3@     ��@      �?                             �H@              �?                               @                                      �?        333333>@fffff��@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @      3@      3@                                      �?      �?       @                                                                      �?      @�����I@�����I@                      �?      �?     �Q@      �?       @               @       @       @       @                       @              @fffff�Q@3333�h�@                                      K@      �?       @      �?                       @       @               @       @      �?        fffff�W@�����ȳ@              �?      �?              M@      �?       @      �?                               @       @       @              �?        �����Y@�����u�@              �?      �?              *@      �?              �?                                                              �?       @������Q@     ��@      �?              �?      �?      @      �?              �?       @               @                       @              �?      @fffff�V@     ({@                                     �C@              �?                               @               @       @              �?       @     `I@�����m�@              �?                      @@      �?              �?                                               @              �?       @     �S@     Ҥ@      �?              �?              @              �?                       @                                                      �?������=@������W@      �?                              K@      �?       @      �?       @       @               @       @       @       @      �?      �?      [@ffff���@                                      &@      �?               @      �?      �?      �?      �?      �?      �?                        �����L4@������n@              �?                       @      �?              �?                       @               @       @              �?       @fffffW@�����φ@      �?              �?              �?      �?                                                                                      �?�����YF@�����YF@              �?                      .@      �?       @      �?                                                              �?      @����̜R@������@                      �?              1@      �?       @                       @                       @       @              �?        ������R@33333��@                                      @              �?                       @                       @       @              �?      �?�����yI@����̬l@      �?      �?      �?      �?     �E@      �?       @      �?               @       @       @       @       @              �?             �[@ffff�O�@                                      �?      �?              �?               @                                                       @33333�R@33333�R@                                      *@      �?              �?                                       @                      �?      @�����yT@������@      �?      �?                     �F@      �?       @      �?                                       @       @              �?        �����yW@    @h�@                                      (@      �?              �?       @                               @              �?      �?      �?�����IU@fffff��@      �?      �?                      @      �?              �?                                                              �?      @������Q@�����9w@      �?                              *@      �?                                               @                              �?      @fffffFI@     �@                      �?              ,@      �?               @      �?      �?      �?      �?      �?      �?       @              @ffffff4@fffffFr@      �?                              @      �?                       @                                                      �?      @33333I@33333d@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     @8@     �@                      �?              "@              �?                               @               @       @              �?       @     `H@33333�{@                      �?              :@      �?                               @               @       @       @              �?       @33333CR@     ��@      �?                              @      �?              �?                       @                                      �?      �?ffffffR@     m@      �?                              8@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@�����p~@              �?      �?               @      �?       @      �?                                               @              �?       @      U@33333+�@                      �?      �?     �N@      �?       @      �?       @       @       @                       @      �?      �?      �?�����,Y@ffff���@      �?      �?      �?      �?     �Q@      �?       @                       @       @       @               @      �?      �?        �����9R@ffff��@                      �?              G@      �?       @      �?               @       @       @       @       @       @      �?      �?�����9[@����L��@      �?              �?              1@      �?              �?                                                              �?        ������Q@33333��@      �?                              @      �?                                       @               @       @      �?      �?      @     �Q@fffff�u@                      �?      �?      "@      �?                               @               @       @              �?      �?      @ffffffP@fffff��@                      �?              &@      �?       @      �?               @                       @       @              �?       @     �Y@fffff�@      �?              �?              P@      �?       @      �?       @       @       @                              �?                �����\V@ffff�<�@                                      J@      �?       @      �?       @       @               @       @       @      �?      �?      �?     �[@3333s�@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?�����i\@33333��@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      �?�����Y4@     �^@                      �?      �?      O@      �?       @      �?               @       @       @       @       @      �?      �?       @33333�[@3333�@      �?                              2@      �?                                       @       @                                      �?������K@fffff��@      �?                              @      �?       @      �?                                                              �?       @������R@�����\}@              �?      �?              A@      �?                                       @       @       @              �?                �����P@�����t�@      �?              �?              I@      �?       @      �?                               @       @       @      �?               @������X@    �ó@      �?                             �P@              �?                                       @                      �?              �?33333s=@�������@                                      �?      �?                                                                                       @33333�F@33333�F@                                      D@      �?       @      �?               @       @               @                      �?        �����YW@�����X�@              �?      �?      �?     �M@      �?       @      �?                       @                       @              �?      �?     0V@ffff��@      �?                      �?     �B@      �?                       @       @               @                       @              �?������N@3333���@              �?      �?              �?      �?              �?                                                              �?       @33333cQ@33333cQ@      �?              �?             �P@      �?       @      �?       @       @       @               @       @      �?              �?�����y[@fffff��@      �?                             �M@      �?                                       @                       @      �?      �?        ����̬N@     {�@      �?                              �?      �?                                                                              �?      @fffff�F@fffff�F@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@33333�A@                                      N@              �?               @               @               @       @       @               @������J@����J�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @     @3@33333�U@      �?              �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������8@33333I�@      �?              �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @ffffff9@fffff�@      �?              �?              D@      �?                               @                                              �?      @33333I@     �@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333s3@     `\@                                      @      �?              �?                               @               @              �?      �?�����YU@fffff�z@      �?                              "@              �?                                               @       @              �?       @33333�F@�����,z@      �?                               @              �?               @                                                              @�����Y=@fffffk@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�4@33333S[@              �?                      ;@      �?       @      �?               @       @                                      �?        ����̜U@����¢@      �?      �?      �?              @              �?               @                                                                ������=@fffff�k@      �?                              P@      �?       @      �?                       @       @       @       @      �?      �?      �?�����)Z@������@              �?                      =@      �?       @               @       @                                              �?        fffffFM@�����ۚ@                                     @P@      �?       @      �?       @       @               @                      �?      �?       @fffffvV@ffff�Զ@      �?                              F@              �?                       @       @               @       @      �?      �?      @������J@����̎�@              �?      �?              �?      �?              �?               @                                              �?      @�����S@�����S@      �?              �?      �?      �?      �?              �?                                                              �?      @�����yQ@�����yQ@                      �?      �?      6@      �?       @      �?                                                              �?        33333�R@fffff<�@      �?                             �J@      �?       @                       @       @       @               @       @      �?        �����yR@    ��@      �?              �?      �?      Q@      �?       @                       @       @       @               @      �?      �?        33333�R@3333�@                      �?      �?      R@              �?               @       @       @       @       @       @       @                �����lP@����Y߱@      �?                              :@      �?              �?                       @       @       @       @              �?       @������X@     ң@                                      >@      �?                       @       @       @       @       @       @      �?                fffffVU@�����ģ@              �?                      "@      �?              �?                                       @                      �?       @fffff6T@33333}�@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����L3@�����L3@                                      (@      �?              �?                       @               @       @              �?       @      X@fffff��@      �?              �?      �?      4@      �?       @      �?               @               @       @                              @333333X@����̊�@                      �?              R@      �?       @      �?               @       @       @       @       @      �?      �?       @     P[@����̭�@      �?              �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?ffffff3@������@                              �?      *@      �?       @      �?               @       @               @       @      �?      �?      �?�����	Z@fffffL�@      �?              �?      �?     �A@      �?              �?               @               @       @              �?      �?       @�����lV@33333��@      �?              �?      �?      6@      �?       @      �?                       @               @                      �?       @     0V@�����t�@                      �?      �?     �Q@      �?       @               @       @       @       @       @               @               @�����,T@3333��@                                       @      �?               @      �?      �?      �?      �?      �?      �?                             �2@33333�J@      �?              �?              R@      �?       @      �?       @       @               @       @       @       @      �?      �?�����|[@fffff��@                                      J@              �?               @       @       @               @       @       @      �?             `M@������@      �?              �?              @@      �?       @      �?                       @                                      �?       @������S@ffff��@              �?                      1@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�4@������t@                      �?      �?     �Q@      �?       @               @       @       @       @       @       @       @                �����yV@3333�Ƹ@                      �?             �O@      �?       @               @       @                       @       @      �?      �?      �?������S@ffff&��@              �?                      @      �?              �?                       @                                               @������R@�����!{@                      �?              R@              �?                       @       @               @       @       @      �?       @�����K@ffff�®@                      �?      �?      M@      �?       @      �?       @       @                               @              �?        �����YW@�����;�@              �?      �?      �?      H@      �?              �?       @               @       @       @       @              �?       @      Z@����̳@                                       @      �?                                                                                      @�����9F@�����w@              �?                      >@      �?       @      �?       @       @       @                                              �?������V@����L��@      �?              �?      �?      M@      �?                               @               @       @       @      �?      �?      �?������R@�����̰@              �?                      G@      �?              �?               @                       @       @      �?              �?     �W@33333H�@      �?              �?      �?     �M@              �?               @               @                              �?              @ffffffA@33333�@      �?      �?                     �B@              �?                       @       @                                               @33333SB@     ��@              �?      �?              @      �?       @      �?                                               @              �?       @fffffU@fffff�}@      �?              �?      �?     �M@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@fffff�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      �?�����4@33333�W@                                      5@      �?              �?               @       @                       @              �?       @33333�V@������@      �?                      �?      �?      �?                               @                                              �?       @33333�H@33333�H@      �?              �?      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�����L9@fffff!�@                                     �G@      �?              �?       @               @       @       @       @      �?      �?       @������Y@�����z�@                                      O@              �?                       @       @                       @       @      �?      �?������E@fffffy�@      �?      �?                      "@      �?       @      �?                                               @              �?       @33333CU@     T�@                      �?      �?     @Q@              �?                       @       @               @       @       @      �?      �?�����yK@     y�@      �?              �?              7@      �?       @      �?       @       @       @               @                      �?       @     �X@������@      �?              �?      �?      R@              �?               @       @       @       @               @       @      �?      �?������K@33333S�@                      �?              L@      �?       @      �?                       @       @       @       @       @                ������Y@����Yp�@      �?              �?      �?      N@      �?                       @       @               @       @       @              �?      �?33333�S@fffff7�@      �?              �?      �?      A@              �?                               @       @       @                      �?       @�����lF@fffff��@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@������I@                                     �G@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @����̌4@�������@      �?              �?      �?      N@      �?                               @               @       @       @       @                �����<S@3333�@                              �?      *@      �?       @               @       @       @       @       @       @       @              �?�����<V@     '�@                                      M@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?33333�8@     ��@                                      &@      �?       @                                                       @              �?      @�����yM@�����̂@                                      .@      �?                       @               @       @                                       @�����yM@33333ٍ@      �?              �?      �?     �D@      �?       @      �?                       @       @       @       @      �?      �?       @fffff�Y@����Yu�@      �?                      �?      6@      �?              �?               @       @               @                      �?       @�����YV@     F�@      �?              �?      �?      ?@      �?       @               @       @               @               @      �?      �?             �R@     Q�@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?                             @4@33333wt@              �?                       @      �?       @      �?                       @                       @              �?       @33333#V@     hf@                                     �I@      �?       @      �?       @       @       @               @       @      �?                ������Z@ffff�0�@                                      @              �?               @                                                      �?      @fffff&=@33333�[@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff3@�����YW@                                      *@      �?       @      �?       @                                                      �?      �?      T@fffff�@                                      @      �?       @      �?                                                              �?       @����̼R@����̌j@              �?                      G@      �?       @      �?       @       @       @               @       @      �?      �?       @     �[@�����
�@                      �?      �?      R@      �?                       @       @       @       @       @       @       @                33333SU@33333�@              �?                      �?      �?       @      �?                                                              �?       @����̌R@����̌R@      �?              �?             �A@      �?       @      �?                               @       @                      �?      �?     �V@3333�H�@                      �?             �P@      �?       @                       @       @       @       @       @       @                ������U@�������@      �?              �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?      �?33333#]@����Lؿ@      �?                              $@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @      8@�����Ql@      �?              �?      �?     �K@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@�����g�@      �?              �?      �?     �C@              �?                                                              �?      �?      �?     @9@     ��@      �?              �?             �O@      �?       @      �?               @       @               @       @              �?       @������Y@����,�@      �?              �?             �G@      �?       @      �?       @               @       @       @       @      �?      �?      �?fffff�[@����̛�@      �?              �?              ,@      �?       @      �?                                       @                      �?       @fffff�U@33333N�@      �?      �?      �?      �?      Q@      �?       @      �?                       @       @       @       @      �?      �?      �?������Z@�����Ӽ@      �?              �?             �N@      �?       @                       @       @               @       @      �?      �?       @33333�S@�����2�@                      �?      �?      M@              �?                               @       @       @       @       @      �?      �?     �K@����̽�@              �?                      @      �?       @      �?                                               @              �?       @fffff&U@������v@      �?                              @      �?              �?                                                              �?       @     pQ@�����It@      �?                              4@      �?       @      �?                       @               @                      �?      �?����̬V@fffff՛@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@����̌?@      �?      �?                      @      �?       @      �?                       @               @                               @33333�V@�����r@                      �?      �?      M@      �?       @      �?               @       @               @       @      �?      �?      �?�����LZ@fffffQ�@              �?      �?      �?      ?@      �?              �?                       @       @       @       @              �?       @������X@�������@              �?      �?      �?      H@              �?                       @                                      �?                fffff�=@     ��@      �?                              @      �?                       @                       @       @                      �?      �?�����P@�����th@                                      (@      �?               @      �?      �?      �?      �?      �?      �?                        33333s3@fffffnl@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?       @                �����Y3@33333c�@      �?              �?      �?      R@      �?       @      �?               @                       @              �?      �?       @�����lV@3333�@      �?      �?                     �I@      �?       @      �?                       @               @       @              �?       @33333sX@����L1�@                              �?      F@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@����� �@      �?                              .@              �?                                       @                              �?       @33333�=@     d{@      �?              �?              R@      �?       @      �?       @       @               @       @       @       @      �?      �?�����<[@     þ@      �?              �?             �Q@      �?       @                       @       @       @       @       @       @              �?�����U@�����D�@              �?                      0@      �?       @               @                                                      �?       @�����K@     ȋ@      �?              �?      �?     �G@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @����̌8@�����!�@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @3333333@3333333@                                      (@      �?       @               @               @       @                              �?      @33333�N@     N�@      �?                              5@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@ffffffx@              �?                      �?      �?                       @               @                                      �?       @fffff�K@fffff�K@                                      �?      �?                                                                                        33333F@33333F@      �?                              O@      �?       @       @      �?      �?      �?      �?      �?      �?       @                ffffff7@�����V�@                      �?      �?     �A@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?ffffff9@fffff��@      �?                              *@      �?       @      �?                               @       @       @              �?      @     �X@�����V�@      �?              �?      �?      O@      �?                       @       @       @       @       @       @       @               @fffff�U@    @_�@                      �?      �?      @      �?       @      �?               @                       @       @              �?       @�����|X@     x@                                      6@              �?                       @                       @       @              �?       @�����,I@fffff+�@      �?                              @      �?              �?                                                              �?       @fffffFQ@     0{@                                      "@      �?       @      �?                                       @       @                       @������W@     ʊ@                      �?              3@      �?       @      �?                       @                       @                      @�����iV@33333��@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?             @9@�����Ĝ@                      �?              $@      �?                                       @               @       @              �?      �?33333�P@33333i�@      �?                              D@      �?                       @               @                       @                       @������P@     V�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?       @������3@������3@      �?                              I@              �?               @       @                                              �?      @     �A@�����ٛ@                      �?              E@      �?       @                                                                      �?       @      I@����L7�@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?       @     �\@3333�t�@                      �?              Q@      �?       @      �?       @       @       @       @       @       @       @                ������\@���̌��@                      �?      �?     �M@      �?       @      �?               @               @               @              �?        �����)X@�����̵@      �?                              D@      �?              �?               @               @               @      �?      �?      �?ffffffV@����L@�@      �?      �?                      :@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����L3@33333�@                      �?      �?      R@      �?              �?       @       @       @       @       @       @       @      �?        �����)[@����Y.�@                                       @      �?              �?                                       @                      �?      @������S@fffffc@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @3333334@3333334@                                     �D@      �?       @      �?               @       @               @       @              �?       @33333�Z@3333s[�@      �?      �?      �?      �?      4@      �?              �?       @               @       @               @      �?              �?33333�W@33333i�@                      �?      �?      9@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@�����`~@      �?                      �?      O@      �?                       @       @                                      �?                33333L@ffff�?�@      �?                      �?      K@      �?              �?       @       @               @       @       @      �?      �?       @fffffvZ@ffff�¶@      �?      �?      �?             �Q@      �?       @      �?       @       @       @       @       @       @       @      �?        33333�\@�����P�@      �?                              �?      �?              �?                                                                      @fffff�Q@fffff�Q@      �?              �?              L@      �?       @      �?       @       @       @                              �?      �?       @�����IW@3333�@                      �?      �?      *@      �?               @      �?      �?      �?      �?      �?      �?       @      �?             �3@fffff�n@      �?                      �?      (@      �?                       @                               @       @              �?      @fffffvQ@     ,�@      �?                              �?      �?       @      �?                       @               @       @              �?       @�����\Y@�����\Y@                      �?      �?      @              �?               @                       @                                      @33333SA@33333�n@      �?              �?      �?      7@      �?              �?       @                       @       @       @              �?       @fffff�X@�����6�@      �?                              2@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@�����y@      �?              �?      �?     �N@      �?                       @       @       @       @                       @      �?        33333Q@    @>�@      �?              �?      �?      @@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?33333s3@fffff�@                      �?              Q@      �?                               @               @       @               @                fffffP@    @�@                      �?              Q@      �?       @      �?               @       @       @                       @              �?����̌V@ffff���@                              �?       @      �?                       @                                       @              �?      �?������N@�����|_@                                      =@      �?       @      �?                                                              �?      �?      S@    �N�@                                      C@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?       @     @8@33333��@      �?      �?      �?              *@      �?              �?                                                                        ����̜Q@����̈�@                      �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?                      @33333s4@     j�@                      �?      �?      J@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?       @ffffff4@�����
�@      �?                      �?      �?      �?                       @                                                              @�����LI@�����LI@      �?              �?      �?      :@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?fffff&3@     �@                      �?      �?      8@      �?                       @                       @                                       @33333�K@fffff��@                                     �A@      �?       @               @               @       @       @       @      �?      �?      �?�����|U@33333L�@      �?      �?                      3@      �?       @      �?       @                               @                      �?       @fffff�V@     �@                      �?              F@      �?       @      �?       @       @       @       @                              �?      �?fffff�W@������@      �?                             �M@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @      9@     ��@                                     �B@              �?                               @                       @              �?      �?�����D@fffff�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����L4@�����L4@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?ffffff8@�������@              �?                      @      �?                               @                                              �?      @fffff�I@�����5z@      �?              �?      �?     �Q@      �?       @      �?       @       @                       @                      �?      �?33333cX@�����@                      �?             �H@      �?       @      �?       @                               @       @              �?      @fffff6Y@����Y�@      �?                               @      �?                       @       @                                              �?      @������J@�����	[@      �?                              @      �?                                                               @                       @fffff&K@�����ih@      �?                              (@      �?       @       @      �?      �?      �?      �?      �?      �?                       @      9@33333�s@                      �?      �?      3@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        fffff�8@33333;}@                                      �?      �?              �?               @                                              �?       @����̬R@����̬R@      �?                      �?     �A@      �?                                               @       @       @      �?      �?      @fffffR@����L~�@      �?                              F@      �?              �?               @               @       @       @                       @33333#Y@ffff&.�@      �?      �?      �?              &@      �?              �?                                                              �?       @����̌Q@������@                                       @      �?                               @                                              �?      �?fffff�H@fffff�V@      �?              �?              $@      �?       @      �?                       @               @       @              �?       @     �X@     7�@                      �?      �?       @      �?              �?                       @               @       @              �?       @����̌W@fffffJ�@      �?              �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff&4@     �d@      �?              �?      �?      N@      �?                       @       @       @                               @                     @N@ffff�ܬ@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      �?������3@33333[a@      �?              �?             �P@      �?              �?       @       @                       @       @      �?      �?      �?�����9Y@ffff&M�@      �?                      �?      9@      �?               @      �?      �?      �?      �?      �?      �?                      @������4@33333�|@      �?              �?      �?      O@      �?               @      �?      �?      �?      �?      �?      �?       @                33333s4@fffffE�@      �?      �?      �?      �?      L@      �?       @      �?       @               @               @       @      �?      �?        33333#Z@ffff���@      �?              �?      �?      $@      �?                                       @               @                              @�����N@     ��@      �?              �?      �?      I@      �?       @      �?       @               @               @       @                      �?�����|Z@�����ݴ@      �?                              @              �?               @               @                              �?              @fffff�A@����̌p@      �?                              6@      �?       @               @       @                                                       @     �M@����̚�@      �?              �?              A@      �?       @      �?               @                               @                      @fffff6V@    �p�@      �?              �?              =@      �?       @      �?               @       @                                      �?       @33333sU@    ��@                      �?      �?     �Q@      �?       @      �?       @       @       @               @               @                      Y@ffff�v�@                                      7@      �?               @      �?      �?      �?      �?      �?      �?              �?        �����L4@�����i}@                      �?              E@      �?               @      �?      �?      �?      �?      �?      �?                      �?�����Y4@33333/�@      �?      �?      �?             �N@      �?       @      �?               @                                              �?       @������T@�����(�@      �?              �?      �?      R@      �?       @      �?       @       @       @       @               @       @              �?������Y@3333�]�@                      �?      �?      *@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?              9@     �t@      �?              �?              Q@      �?       @      �?       @       @               @       @       @              �?       @������Z@ffff昼@      �?              �?             �Q@      �?       @      �?               @               @       @       @       @      �?      �?�����	Z@����Lż@                      �?      �?      $@      �?              �?                                       @       @              �?       @fffff6V@������@                      �?      �?     @P@      �?       @      �?       @               @       @       @       @       @               @33333S[@���̌��@                      �?              G@      �?       @               @                                                               @����̌J@�����7�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @33333s3@     PQ@      �?              �?              @      �?       @      �?               @                       @       @              �?       @�����Y@33333Cz@                      �?              $@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@�����g@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�2@�����lt@                      �?      �?      1@      �?                       @                       @                              �?      �?����̬K@     Č@                                      �?      �?                                       @                                      �?      @�����9I@�����9I@                                      G@      �?       @               @               @               @       @       @              @������S@������@                      �?      �?      R@      �?       @      �?       @       @                       @               @      �?        ������W@ffff&*�@                      �?             �C@      �?              �?       @               @       @       @       @      �?      �?      �?�����,Z@�����&�@      �?                              �?      �?                                                                                       @      F@      F@                              �?      O@      �?       @      �?                       @               @       @      �?      �?       @�����	Y@ffff��@                                      �?      �?                                                               @              �?       @      L@      L@      �?                              &@      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@     �j@                      �?      �?      &@      �?       @                                       @               @              �?       @fffff�P@fffff&�@      �?                              2@              �?                       @       @                                      �?      �?     �@@     ��@      �?      �?                      6@      �?       @      �?                                       @       @              �?       @�����,X@ffff�E�@                                      @      �?       @                                       @       @                               @fffff&P@fffff�e@      �?              �?      �?      @              �?               @                       @                              �?       @     @A@     tq@      �?      �?      �?      �?     �P@      �?       @               @       @       @       @       @               @              �?������S@�����"�@      �?      �?                     �G@      �?              �?       @                                       @                      @     `U@�������@                                      R@      �?              �?       @       @       @       @       @       @       @      �?       @�����y[@33333Ƚ@                      �?      �?      R@      �?              �?       @       @       @       @       @       @       @      �?      �?     `[@ffff殾@                      �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @                ����̌3@�����ݖ@                                     �N@      �?       @      �?       @       @       @       @       @       @      �?      �?      @fffff�\@ffff�Q�@      �?              �?              ,@      �?       @                                       @       @                      �?      �?fffff�P@     ��@      �?                      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@fffff�p@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                       @33333s3@33333s3@                      �?      �?      @      �?       @                                                                              @�����lI@������m@      �?      �?      �?              @      �?       @      �?                                                              �?       @fffff�R@     T~@      �?                              A@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����:@����̢�@      �?                              �?      �?                                                                              �?      @�����yF@�����yF@                                      (@      �?                               @               @                              �?       @fffff&K@     t�@                      �?      �?      1@      �?       @      �?       @               @               @       @              �?       @�����Z@     >�@                                      @      �?                                       @       @               @                        ffffffO@�����$z@                      �?      �?      @              �?                       @                                              �?       @     �>@fffff�d@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333s4@33333s4@      �?                              7@      �?       @      �?                       @       @       @       @              �?      @33333Z@33333L�@                      �?      �?      4@      �?       @       @      �?      �?      �?      �?      �?      �?              �?        ����̌9@fffff�@                      �?      �?      R@      �?       @      �?       @       @               @                       @      �?        fffff�V@fffff��@                                      @      �?       @      �?                                                                       @fffff�R@�����!u@              �?      �?              ;@      �?              �?       @                                                      �?        ������R@fffff%�@      �?      �?                       @      �?              �?       @                       @       @       @                      �?33333Y@������@      �?              �?             �Q@      �?       @      �?       @       @               @                       @      �?      �?      V@3333sb�@              �?                      @      �?                               @       @               @                      �?       @�����<P@fffff�~@      �?                             �M@      �?       @      �?               @       @       @       @       @              �?       @fffff�[@    �w�@      �?              �?      �?     �J@      �?       @               @                       @               @                       @fffff�Q@������@                      �?      �?      0@      �?              �?       @               @               @       @                        �����,Y@�����ʗ@                                       @      �?       @      �?                                                              �?       @33333�R@������d@      �?              �?              ,@      �?                                               @                                        ffffffH@33333Ä@                                      B@      �?       @                               @                              �?               @fffff�K@     V�@                      �?      �?     �P@      �?       @               @       @       @       @       @       @       @              �?�����yV@�����F�@                                     �P@              �?                               @       @       @       @              �?      �?33333�J@����L��@      �?              �?      �?      R@      �?       @               @                                               @                fffff�K@33333�@      �?                              I@      �?       @       @      �?      �?      �?      �?      �?      �?       @                fffff�8@     ��@                      �?      �?      *@      �?                       @               @                       @              �?      @33333�O@fffff��@                                       @      �?                                                                              �?      @������F@ffffffZ@                      �?      �?     �D@      �?               @      �?      �?      �?      �?      �?      �?       @                �����L3@33333#�@      �?      �?      �?              �?      �?              �?                                                                      @fffff�Q@fffff�Q@      �?              �?              @      �?              �?                                                              �?       @33333�Q@33333j@              �?                     �B@      �?       @      �?       @       @                       @       @              �?             �Z@    ���@                      �?              I@      �?       @      �?       @               @               @       @      �?      �?      @�����Z@ffff�p�@      �?                      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�3@fffffԓ@                      �?             �J@      �?       @      �?               @       @       @       @       @      �?      �?        33333�[@    ���@      �?                              I@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?fffff&4@fffff�@                                      &@      �?                                               @       @       @                      @     �Q@fffff�@      �?      �?                      P@      �?       @      �?                       @       @       @       @      �?               @fffff�Y@���� �@                      �?              L@      �?              �?                       @       @       @       @              �?       @����̬X@    �%�@                      �?      �?      K@      �?       @      �?       @       @                       @       @              �?        fffffZ@������@      �?                              2@              �?               @               @                                              @������@@�����2�@      �?                      �?      �?              �?                                                                               @     �8@     �8@      �?              �?      �?      I@      �?              �?               @       @       @       @       @      �?      �?        ������Y@ffffft�@      �?                              @      �?                                                       @                              @33333�K@������c@      �?              �?      �?      @      �?                                                                                       @ffffffF@�����4e@      �?                               @      �?                                                                                        33333sF@33333�[@      �?                      �?     �A@      �?              �?                       @               @              �?      �?       @�����IU@33333��@                                      "@      �?               @      �?      �?      �?      �?      �?      �?                      @�����3@����̴c@      �?                      �?      @      �?                       @                                                      �?       @33333�H@�����g@                      �?      �?      ;@      �?              �?       @                                                              @������R@fffffў@                                      &@      �?       @      �?                                                              �?       @      S@�����/�@      �?              �?      �?       @      �?                                                                      �?      �?      @������E@     �u@      �?                              2@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @     �7@     �z@                      �?      �?     �D@      �?                               @               @               @      �?      �?             �P@33333Q�@                              �?      0@      �?       @      �?                               @                      �?      �?      �?     �S@�������@                                      �?              �?                                                                      �?      @fffff�8@fffff�8@      �?                              &@      �?              �?               @                                              �?      @������R@33333�@                      �?      �?     �K@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����L4@33333ܐ@      �?              �?      �?     �O@      �?       @      �?               @                               @      �?      �?       @fffff�V@3333���@                              �?     �I@              �?               @               @       @       @       @      �?                33333N@     
�@                      �?      �?      �?      �?                                                                              �?        �����,F@�����,F@                                      �?      �?       @                                                                      �?       @�����I@�����I@      �?                             �P@      �?                       @       @                                      �?      �?      @ffffffK@fffff�@                      �?      �?      J@      �?              �?               @       @       @                                        33333sU@����LQ�@      �?              �?      �?     @P@      �?       @                       @       @       @       @       @       @      �?        �����U@    �̴@              �?      �?              @      �?              �?                                       @                      �?       @�����T@�����l@                      �?      �?      2@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?fffff�8@�����u}@                                      ;@      �?                       @       @                                              �?      @�����YL@�����ә@      �?                               @      �?                                                                              �?      �?      G@      U@                                      E@      �?                       @       @       @       @               @      �?              �?�����yR@������@      �?              �?      �?      8@      �?                       @               @                              �?      �?      �?      L@     ��@                      �?              L@      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @�����L8@����̶�@      �?              �?      �?      I@      �?       @                               @                              �?                33333sK@33333l�@      �?      �?      �?             �M@              �?                       @                       @       @              �?       @      I@ffff�j�@      �?              �?              =@              �?                                               @       @              �?       @33333�F@�����є@      �?                              :@      �?              �?               @                                      �?                     �R@fffff��@                      �?             �Q@      �?       @               @       @       @       @       @       @       @                ������U@����Yݸ@                                      0@      �?       @                                                       @              �?        fffff�O@33333��@      �?                              Q@      �?       @               @       @       @                       @      �?              �?     0S@    @q�@      �?              �?              8@      �?              �?       @                       @               @              �?       @     PV@fffffD�@      �?      �?      �?      �?      8@      �?       @      �?       @                                                      �?       @fffff�S@     �@                                      A@      �?              �?               @                                              �?      �?�����|R@ffff渣@      �?                              D@      �?                       @       @               @                              �?      @33333�N@33333��@      �?              �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @ffffff9@33333؛@                      �?      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?       @                     �3@33333��@                                      6@              �?                               @               @       @              �?       @�����LI@33333Ő@              �?      �?              (@      �?                       @               @       @       @       @      �?      �?       @������S@�����~�@                      �?             �G@      �?              �?                       @                       @              �?       @33333SU@����L��@                                       @      �?                       @                               @       @              �?       @     �Q@�����\b@      �?              �?      �?      6@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@     {@      �?      �?                      $@      �?              �?               @                                              �?       @fffff6R@33333��@                      �?      �?      @      �?                                                                                      @     �F@33333�q@      �?                              @      �?       @      �?                               @               @              �?        ������U@�����R�@      �?              �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����8@������@      �?              �?      �?      F@              �?                               @       @       @       @      �?      �?       @fffff&K@33333�@      �?      �?                      9@      �?       @      �?               @                       @                      �?       @�����<V@fffff�@      �?              �?      �?     �D@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @      4@fffff~�@                                      �?      �?              �?                                                              �?       @fffff�Q@fffff�Q@              �?                      �?      �?              �?                                                              �?       @������Q@������Q@      �?                              6@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����L4@������}@      �?              �?      �?      D@              �?                       @       @       @       @       @      �?              @fffff&N@     !�@      �?      �?      �?              >@      �?              �?               @       @                                      �?      @������S@����Lz�@      �?              �?             �L@      �?                       @       @               @                       @      �?       @     �M@����L��@              �?                      N@      �?       @      �?       @                               @       @      �?      �?        �����YY@����� �@                      �?      �?      2@      �?                                                       @                              @������K@33333�@      �?                      �?     �D@      �?                       @       @       @               @              �?              @����̌Q@������@      �?                              �?      �?                                                               @                      @fffff�K@fffff�K@      �?                              ;@      �?       @                                                                              @     �H@fffff-�@      �?              �?      �?     �P@              �?                               @       @       @       @       @                33333SK@     `�@      �?      �?                     �L@      �?       @      �?       @                       @               @       @               @     pW@���̌��@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@     �K@                                      P@      �?       @      �?                       @               @       @      �?      �?      �?33333Y@33333n�@      �?      �?                      >@      �?                       @       @                       @       @              �?       @     �R@�����~�@                                      4@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�����Y3@     {@                                      0@      �?                       @                                                      �?       @33333I@     ҇@      �?                              �?              �?                                       @                                      @fffff&=@fffff&=@      �?              �?      �?     @P@      �?       @               @       @                               @       @      �?      @33333cQ@ffff&k�@                                      $@      �?       @      �?                                                              �?      @     �R@fffffJ�@                      �?      �?      5@              �?               @               @               @       @      �?      �?       @������K@33333�@      �?                              �?      �?              �?                                                                       @�����|Q@�����|Q@                      �?              7@      �?                                               @       @              �?                      N@������@                      �?      �?      O@      �?                       @               @                              �?              �?     `K@3333�ª@                      �?      �?     �P@      �?       @      �?               @       @       @       @       @      �?      �?      �?fffff\@3333sܼ@                                     �@@      �?       @               @                       @                      �?               @33333�M@33333��@      �?              �?              R@      �?       @      �?               @       @       @       @       @       @      �?       @�����[@    �'�@      �?      �?      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        ����̼\@33333�@                      �?      �?      &@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @      4@33333�h@      �?              �?              R@      �?       @               @       @       @       @       @       @       @      �?      �?     �V@3333s�@      �?              �?             �Q@      �?              �?       @       @       @       @       @       @      �?      �?             `[@ffff�n�@                      �?      �?     �@@      �?                       @       @       @                              �?      �?      @�����9M@�������@      �?      �?      �?             �L@      �?       @      �?               @       @                       @              �?             �W@����3�@      �?              �?              L@      �?       @      �?       @                               @       @      �?      �?       @33333#Y@3333�@                                      *@      �?              �?               @       @                                      �?       @�����IT@fffff@      �?      �?                      .@      �?       @      �?                                                                       @������R@������@                                      *@      �?              �?               @       @                                      �?       @     �S@�����^�@                                      �?      �?              �?                                                                       @�����)Q@�����)Q@      �?                              6@      �?       @      �?       @                               @       @              �?        fffffVY@33333�@                                      D@      �?              �?               @                                                      �?33333�R@fffff7�@      �?      �?      �?              G@              �?                       @       @       @       @       @      �?      �?        33333�M@����L�@      �?              �?      �?      >@      �?               @      �?      �?      �?      �?      �?      �?       @              @     @5@33333?�@      �?                              "@      �?              �?                               @       @       @              �?        ������W@�����ۉ@              �?      �?             �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����4@33333��@      �?              �?      �?      2@      �?              �?                               @               @              �?       @ffffffU@     �@      �?              �?      �?      R@      �?              �?       @       @               @       @       @       @                     `Z@���̌��@                      �?      �?      .@      �?                               @       @       @       @       @                              S@fffff�@      �?              �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @              �?ffffff3@     M�@      �?              �?      �?     �N@      �?               @      �?      �?      �?      �?      �?      �?       @              �?����̌4@�����g�@                      �?              R@      �?       @      �?               @       @       @       @       @      �?      �?              [@�����C�@                                      >@      �?                       @       @                                              �?        fffff�K@fffff�@      �?                             �H@      �?       @      �?               @               @       @       @      �?      �?        ������Z@����0�@                      �?               @      �?              �?       @                       @                              �?       @�����	T@�����Qh@                                      @      �?       @      �?                                                              �?      �?fffff�R@33333�p@      �?              �?      �?     �H@      �?       @      �?                       @               @       @              �?       @33333�X@3333s�@                                      ,@      �?              �?                                                              �?      �?     �Q@     ��@                                      C@      �?       @      �?                       @       @       @       @              �?       @������Y@     )�@      �?                              R@      �?       @               @       @       @       @       @       @       @                ������U@�����P�@              �?      �?              R@      �?       @      �?       @       @                       @       @      �?      �?        fffff�Z@fffff��@      �?                              �?      �?       @      �?                                                              �?       @fffff�R@fffff�R@      �?              �?      �?      P@      �?       @      �?               @       @       @       @       @       @      �?      �?�����L[@ffff&U�@      �?              �?      �?      $@      �?                               @                                      �?              @fffff�H@33333�}@                              �?      (@      �?       @      �?                                                              �?       @fffff&S@     �@                              �?      (@      �?       @      �?               @       @               @       @              �?       @33333SZ@������@                      �?      �?      J@      �?              �?       @               @               @       @      �?               @33333Y@3333s|�@              �?                      L@      �?       @      �?               @       @               @       @      �?      �?             0Z@ffff���@                      �?      �?     �M@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @33333s9@33333��@                                     �C@      �?                               @                       @              �?      �?      �?�����LM@     a�@      �?                              �?      �?                                                                              �?        ����̌F@����̌F@      �?      �?                       @      �?              �?               @                                              �?       @����̬R@����̬d@                                       @      �?       @                                       @                              �?      @�����,K@33333C]@                                      @      �?               @      �?      �?      �?      �?      �?      �?                        33333�4@     `U@      �?              �?             �P@      �?       @      �?               @       @                       @      �?               @33333�W@fffff��@                      �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?�����Y4@�������@      �?              �?             �L@      �?       @      �?       @       @       @       @       @                      �?       @33333�Y@    �%�@      �?              �?      �?      @@      �?       @      �?       @                               @       @              �?      �?33333�X@����L	�@      �?              �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @     �3@     �@              �?      �?              @      �?              �?                               @       @                      �?      @������T@fffff�p@      �?                             �D@      �?              �?               @               @       @       @       @      �?      �?������X@����Y|�@      �?              �?              ?@      �?                                       @       @               @              �?      �?������P@33333��@      �?      �?      �?              Q@      �?       @      �?                       @                                      �?      �?fffffT@����Lյ@              �?                      �?      �?              �?                                       @                      �?       @������S@������S@      �?              �?              "@      �?                       @       @               @       @                      �?      @�����<Q@����̎�@                      �?      �?      Q@      �?       @               @       @       @       @               @      �?      �?       @����̜S@����Yմ@              �?      �?             �Q@      �?              �?               @       @               @       @       @      �?       @������X@    �-�@      �?              �?      �?      A@      �?              �?                       @               @                      �?      @33333U@ffff滦@                                      8@      �?                       @                       @                                      �?�����,L@����̔�@                                      H@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?�����9@     N�@                                      @      �?       @      �?                                                                      @������R@     ~@                      �?              A@      �?       @       @      �?      �?      �?      �?      �?      �?                       @33333�8@�����a�@                              �?      �?      �?                                                                                      @������F@������F@                      �?              P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @����̌9@�����˚@      �?      �?                      I@      �?       @      �?                                       @       @              �?       @������W@3333�в@      �?      �?      �?             �Q@      �?       @      �?       @       @       @       @                      �?      �?       @      W@33333��@                      �?             @P@      �?       @      �?       @               @               @       @              �?       @33333CZ@3333��@                                      4@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@33333oy@      �?              �?             �O@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        33333�3@33333K�@      �?              �?              >@      �?                                       @                                      �?      @      I@������@                                     �B@              �?                                       @                                      �?������<@fffffl�@                      �?      �?     �L@      �?       @      �?               @                       @       @              �?       @fffff&Y@3333��@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @ffffff3@ffffff3@      �?              �?      �?      �?      �?       @      �?                                                              �?       @     �R@     �R@              �?                       @      �?       @      �?               @                               @                       @     `V@     0d@      �?                              L@      �?       @      �?       @       @                                              �?       @������U@fffff:�@      �?              �?              �?      �?              �?                               @       @                      �?       @333333U@333333U@                                      "@      �?               @      �?      �?      �?      �?      �?      �?              �?       @     �3@33333[f@      �?                      �?      (@      �?               @      �?      �?      �?      �?      �?      �?                      �?�����5@�����ym@      �?      �?      �?              8@              �?               @                                       @                        ����̌C@fffffZ�@      �?                              1@      �?              �?                       @                                      �?       @�����)S@33333��@      �?                              @      �?              �?                       @               @       @                              X@������~@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      �?33333�3@33333�3@      �?                             �I@      �?       @               @       @       @       @       @              �?      �?      �?�����IT@33333�@      �?                      �?      5@      �?       @       @      �?      �?      �?      �?      �?      �?                      @33333�8@fffff2}@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                        3333334@3333334@      �?                              �?      �?       @      �?                                       @                      �?      @�����)U@�����)U@                              �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?����̌4@33333�L@      �?                              (@      �?       @      �?                       @               @                      �?       @33333cV@     �@                      �?              9@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        3333334@fffff�@                      �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����8@     ��@              �?      �?              R@      �?       @      �?               @       @               @       @      �?      �?      �?     pZ@�����ͽ@                      �?      �?      4@      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����`y@                      �?      �?     �F@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?fffff�8@33333M�@      �?                      �?       @      �?               @      �?      �?      �?      �?      �?      �?                      @     @3@�����,H@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                3333339@fffff�@                                      (@      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@������p@                                     �G@      �?       @               @       @               @               @       @              @33333�R@�����P�@      �?                              ?@      �?       @      �?               @       @               @       @      �?      �?       @������Y@ffff���@                                      .@      �?              �?               @                       @                      �?        ������T@     ��@      �?                              �?      �?                       @                                                               @������G@������G@      �?              �?      �?     �P@      �?                       @       @       @       @       @              �?      �?       @fffff�R@     ��@      �?                              (@      �?       @                               @               @       @                             �R@fffff؉@                                      K@      �?       @      �?               @                       @       @       @      �?        �����LX@3333s	�@                      �?      �?     �C@      �?       @      �?               @       @       @                      �?      �?       @33333cV@ffff�$�@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @�����L4@������D@                              �?      :@              �?                               @                                      �?      @������=@     ��@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?fffff&\@ffff���@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�3@fffffQ@      �?      �?      �?      �?      M@      �?       @      �?       @       @               @                      �?      �?        fffffvV@    ��@      �?                      �?      �?      �?              �?                                       @       @              �?       @fffff�V@fffff�V@      �?                      �?      7@              �?               @       @               @                      �?                33333SD@33333��@      �?                      �?      �?      �?                       @       @               @               @              �?        ����̜Q@����̜Q@                      �?              Q@      �?       @      �?                       @               @               @      �?        �����|V@����LV�@                                      @@      �?               @      �?      �?      �?      �?      �?      �?                        fffff�3@fffff̂@                                      @      �?                                                                                      @33333�F@������g@                              �?     �E@      �?                       @       @                               @              �?       @������O@����b�@      �?              �?             �A@      �?       @      �?                                                              �?       @������R@fffff �@      �?              �?              R@      �?       @      �?       @               @       @       @       @       @      �?      �?������[@����l�@      �?              �?      �?      �?              �?                       @                                                       @333333>@333333>@      �?      �?      �?      �?     �G@      �?              �?               @                       @              �?      �?        �����<U@����d�@      �?              �?      �?      I@      �?                       @                       @       @       @      �?               @     �R@33333s�@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      �?fffff&4@fffff&4@      �?                              >@      �?       @               @                                       @              �?      @      P@����́�@      �?                              @              �?               @               @       @                                      @      D@fffff�k@                      �?              E@      �?       @               @               @       @       @       @       @              �?fffffU@33333�@              �?                     �A@      �?       @      �?       @       @       @               @       @      �?      �?       @fffff[@����L�@                      �?      �?      0@      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y3@fffff>q@                                     �G@              �?               @       @               @                      �?              �?33333�C@������@                                      @      �?                       @       @       @                                               @33333�N@fffffn{@                      �?      �?      $@      �?       @      �?                                               @                       @�����|U@�����Ԋ@                                      2@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@�����py@                                      >@      �?       @      �?               @       @       @       @       @      �?              �?����̜[@������@      �?              �?             �L@      �?                       @                       @                                       @������K@33333Ǩ@                      �?              @      �?                       @       @                                                      @�����YK@�����am@      �?              �?              I@      �?               @      �?      �?      �?      �?      �?      �?       @               @������3@�������@                      �?              �?      �?                       @       @                                              �?      @fffff�J@fffff�J@      �?              �?             �J@      �?              �?               @                       @       @      �?      �?             �W@3333��@      �?                              (@      �?                                               @       @              �?      �?       @fffff�M@fffff��@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�3@     �F@                              �?       @              �?               @                                       @              �?       @     @C@����̬t@      �?              �?              D@      �?       @      �?               @       @               @       @      �?      �?             �Z@ffff�R�@                                      *@              �?               @                                                      �?        ������>@������x@      �?              �?              &@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����̌4@fffffg@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@������f@                                      �?      �?              �?                                                              �?       @     �Q@     �Q@                      �?      �?      G@      �?              �?                       @       @               @      �?                ����̼V@�������@              �?                      �?              �?                                                                      �?      @������9@������9@                      �?              0@      �?       @      �?               @                       @       @              �?       @      Y@     ��@      �?              �?              @      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @�����9@     `e@      �?              �?             @Q@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@�����M�@                      �?      �?      J@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����7@fffff��@                      �?      �?      �?      �?       @      �?       @               @               @       @              �?       @����̜Y@����̜Y@      �?              �?              ?@      �?                       @       @       @       @               @      �?      �?      �?     �R@ffff��@      �?                             �A@      �?                                                       @                              @     �K@33333j�@                                      A@      �?       @               @       @               @                      �?      �?      @�����P@    �Q�@      �?      �?      �?             �J@      �?       @               @                       @                      �?      �?       @fffffN@����L;�@      �?              �?      �?      A@      �?       @                               @               @       @      �?                �����LS@�������@                                      �?      �?              �?                       @                                               @fffffS@fffffS@              �?                       @      �?              �?                                                              �?       @fffff�Q@�����aa@      �?              �?      �?      I@      �?       @      �?       @       @       @               @       @      �?      �?       @     [@fffff7�@              �?                      I@      �?       @      �?                       @       @       @       @              �?       @�����<Z@����Yf�@      �?                      �?      B@      �?              �?               @                       @       @              �?       @����̬W@     q�@                                      @      �?       @      �?               @                       @                      �?       @     pV@33333E�@                      �?              M@      �?       @      �?       @       @               @       @       @       @      �?      �?fffffF[@ffff���@                                      ?@      �?       @      �?       @       @                       @       @                       @fffffZ@33333�@                                       @      �?                                                                                       @fffff�F@�����U@      �?                               @      �?              �?       @                                                      �?       @������R@fffff�g@      �?              �?      �?      3@      �?       @      �?                               @       @       @      �?      �?       @�����<Y@33333N�@      �?                              @      �?       @      �?               @                               @              �?       @33333�V@�����w@                                      &@      �?                       @                       @                      �?      �?      @�����LK@�����N�@      �?                              �?      �?                                                               @              �?      @������K@������K@                      �?      �?     �Q@      �?       @      �?       @       @       @               @       @       @      �?             @[@������@              �?      �?      �?      8@      �?              �?                       @               @       @       @      �?       @33333#X@ffff殡@      �?                              &@      �?               @      �?      �?      �?      �?      �?      �?       @              �?����̌3@������k@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@33333�a@                      �?      �?      @              �?                       @                               @                      @fffff&D@      W@                                      �?      �?                                                                                      @������E@������E@      �?              �?              @      �?       @      �?               @                                              �?       @     �S@������y@                      �?             �K@      �?       @      �?                       @                                      �?       @     pS@ffff&j�@      �?                             @P@      �?       @      �?       @               @       @       @       @      �?      �?      �?     �[@ffff��@      �?              �?              5@      �?                                                       @                                �����LK@����̔�@      �?                              �?      �?              �?                                                                       @������Q@������Q@      �?              �?      �?      8@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      �?������4@fffffZ}@      �?              �?      �?      9@      �?                               @       @                              �?              @33333�J@�����-�@                      �?      �?      (@              �?                       @                                                      @333333=@�����Qs@      �?                              2@              �?                                                                              @fffff&9@������}@      �?                      �?      ;@      �?       @      �?                               @                              �?       @     �S@����	�@      �?                              $@              �?                               @                                              @     �=@     �o@      �?              �?              $@      �?       @      �?                                       @                      �?       @ffffffU@�����n�@      �?      �?                      F@      �?              �?                       @                                               @fffffvR@�����d�@      �?      �?                      @              �?                               @       @       @                              �?33333�F@     �j@                      �?      �?      <@      �?       @      �?                               @               @      �?      �?       @����̜V@    ���@                                      *@              �?                                                       @              �?       @����̌A@������{@              �?      �?              9@      �?       @               @                       @       @                      �?      �?     `Q@�����b�@      �?              �?      �?      5@      �?       @               @                               @       @      �?      �?        ������R@     7�@                      �?             �N@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     @4@33333��@                      �?             �M@      �?       @      �?                       @       @       @                               @fffffVW@    �
�@      �?              �?               @      �?               @      �?      �?      �?      �?      �?      �?              �?        ����̌3@�����$d@      �?                              $@      �?       @                                               @       @              �?      �?�����	R@     ҈@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                fffff�9@     |�@                                      (@      �?                               @                                              �?       @33333�H@33333�@                      �?      �?      7@      �?              �?       @       @               @                                      @�����U@fffffC�@      �?      �?      �?      �?     �P@      �?       @      �?       @       @       @       @       @       @      �?      �?       @     ]@    @��@      �?      �?      �?             �Q@      �?       @      �?               @       @               @       @              �?       @����̼Y@    ���@      �?              �?      �?      >@      �?       @               @                                                      �?        �����9K@�����Ҙ@                                      B@      �?                       @       @       @       @               @      �?      �?      @33333�R@����L�@      �?                               @      �?              �?                                       @                      �?       @������S@fffff�e@      �?              �?             �@@      �?       @               @       @       @               @                      �?             0R@ffff��@      �?              �?              N@              �?                       @       @       @       @       @              �?        �����N@�������@      �?                              �?      �?       @      �?                                                              �?      @     �R@     �R@      �?                      �?      >@      �?                               @       @               @              �?              �?      P@�����'�@      �?                              K@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�3@�������@                      �?              @      �?                       @               @       @       @       @                             PT@����� �@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?       @     @4@������N@                      �?              &@      �?       @      �?                       @               @       @              �?       @     �X@����̃�@      �?                              N@      �?       @      �?       @       @       @       @       @       @      �?      �?      �?fffff&]@    ���@      �?                              :@      �?              �?               @       @               @                               @33333sV@�����>�@      �?      �?      �?               @              �?                       @       @                       @              �?      @����̬E@fffff6w@                      �?      �?      2@      �?                       @       @               @                      �?      �?      @     �N@�������@                      �?              G@      �?                               @                       @       @              �?      �?fffffFQ@     ��@                              �?      6@              �?                               @               @       @      �?      �?      �?������H@������@      �?                              (@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����4@     �p@      �?      �?                      9@      �?       @      �?               @       @               @       @                      @�����|Z@    ���@                                      $@      �?                               @               @               @      �?              @�����9P@fffffl�@      �?                              =@      �?              �?                       @       @       @       @              �?      �?33333�X@33333�@                                      $@      �?                               @                                                       @������I@     $@      �?              �?      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �3@�����Us@      �?              �?             �M@      �?       @      �?       @       @       @       @       @       @       @               @     p\@    @��@              �?                     �F@      �?       @      �?                       @               @       @      �?      �?        �����	Y@�����k�@                                      B@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?             @3@fffff>�@      �?      �?      �?              M@      �?       @      �?               @                       @       @              �?       @������X@3333���@                      �?      �?      *@      �?                       @                       @                      �?                33333K@fffff�@      �?                      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?�����L9@33333'�@      �?      �?      �?              R@      �?       @                               @               @       @       @      �?      �?�����\R@     Ѵ@      �?                      �?      �?              �?                                                                      �?       @33333�8@33333�8@                                      9@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     �8@����̠�@      �?              �?      �?      1@      �?       @                       @       @       @                              �?      @����̬P@33333Ԑ@                      �?      �?     �Q@              �?                       @       @       @       @       @      �?      �?        333333M@ffff&�@      �?                             �I@      �?       @      �?                       @                                              �?      T@����Y��@      �?              �?              R@      �?               @      �?      �?      �?      �?      �?      �?       @                33333�4@fffffP�@                                      Q@      �?       @               @                                                              @�����9K@    �Ϭ@      �?              �?      �?     �M@      �?       @      �?       @       @               @       @       @       @      �?      @fffff�[@33333��@      �?                              N@      �?                       @       @       @                               @               @33333�N@    �l�@      �?                      �?      "@      �?                                                       @                               @����̬K@     |@                                      "@      �?                       @       @                       @       @              �?       @������R@fffff��@              �?                      L@      �?       @      �?               @       @               @       @                       @     0Z@����YѶ@                      �?              6@      �?                               @       @                                      �?      @�����YK@     k�@                                      H@      �?       @                       @       @       @       @              �?      �?        fffffvR@�������@      �?                              @      �?                                                                              �?      �?ffffffF@ffffff@              �?      �?      �?      ,@      �?       @      �?                                       @       @              �?       @33333�W@33333	�@                                      9@              �?               @       @       @               @       @      �?               @fffff�N@������@                                      N@              �?               @               @                       @      �?      �?       @�����9F@����̫�@                                      @@      �?               @      �?      �?      �?      �?      �?      �?      �?                     �3@33333��@      �?                              8@      �?       @      �?                                       @       @              �?       @fffff�W@3333�%�@                      �?      �?       @              �?                                                                      �?      @ffffff8@fffffFB@      �?                              @      �?       @      �?       @                               @                               @������V@33333�v@                                      @@      �?       @                       @                                              �?       @�����K@fffff.�@      �?                             �C@      �?       @      �?       @       @                       @       @              �?       @������Z@����L��@      �?              �?             �Q@      �?       @      �?       @       @       @               @               @      �?      �?fffff�X@    � �@      �?      �?                      K@      �?       @      �?               @                               @              �?       @33333�V@�����C�@                                      :@      �?                               @       @                                      �?      �?     `K@�������@      �?                              O@      �?       @      �?       @       @                               @      �?      �?        33333W@3333sc�@      �?                              6@      �?       @      �?                                       @       @              �?      �?������W@����q�@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @3333334@     �T@                      �?      �?      6@      �?                       @       @       @                                              @33333�N@333338�@              �?                       @      �?       @      �?                                               @                       @�����LU@     ��@      �?                              "@      �?                       @                       @               @                      @�����<P@fffff�@                      �?      �?     �P@      �?       @      �?       @               @       @       @       @       @      �?      �?     0[@33333��@                                      �?              �?                                                                                     @9@     @9@                      �?             �M@      �?       @      �?       @       @       @       @               @      �?      �?      �?     �Z@����L�@                                     �O@      �?       @      �?               @                       @       @       @                �����\X@     m�@                                      K@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @     �4@�����.�@      �?                      �?      @@      �?       @                       @       @       @       @       @      �?              �?������T@�������@      �?                              �?      �?                               @                                                       @ffffffI@ffffffI@                      �?      �?     �Q@      �?       @               @                       @       @       @       @      �?        fffff&T@33333T�@                      �?      �?      1@      �?       @      �?                                               @              �?       @�����\U@fffff��@      �?                              :@      �?                       @                       @       @       @      �?                     �R@fffffѝ@      �?                              O@      �?       @      �?       @       @       @                                                ����̬V@3333sҵ@                      �?             �E@              �?               @                       @                                              A@fffff��@      �?                              @      �?       @      �?                                               @              �?       @33333�U@�����b�@                                      .@      �?       @      �?               @                       @       @              �?       @�����	Y@     �@                                       @      �?              �?       @               @                                      �?       @�����T@33333#a@                                      �?      �?                                                                                      @fffff�F@fffff�F@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?             �]@����9��@                      �?      �?      M@      �?              �?       @       @                       @       @      �?              �?     �X@ffff�ֶ@                                      =@      �?       @                                               @       @      �?      �?      �?     �Q@33333@�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      �?     �4@     �4@              �?                     �B@      �?       @      �?                                       @       @              �?       @33333#X@�������@                      �?      �?      O@              �?               @       @               @       @               @                �����YH@������@              �?      �?             �Q@      �?              �?       @       @       @       @       @       @       @      �?        �����l[@    @�@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @�����L3@333333F@      �?                               @      �?       @                                               @                      �?       @     �M@�����I{@                                      2@      �?       @      �?               @                       @                      �?      �?     �V@fffffݗ@                                      @      �?              �?               @               @               @              �?       @fffffVV@33333�|@                                      �?      �?                                                                              �?       @�����F@�����F@      �?                              (@      �?                                                                              �?        33333�F@333337�@                                      >@      �?                       @       @       @       @       @              �?              �?������R@33333	�@                                     �F@      �?       @      �?       @       @                               @      �?                     0X@    �Z�@                      �?               @      �?              �?       @       @                       @                               @fffff�V@     �g@                                      "@      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@�����Dg@                                      <@      �?                               @               @                                        33333SK@     ��@                                      A@      �?       @                                       @       @                              @     @P@     ۠@      �?                              @      �?       @       @      �?      �?      �?      �?      �?      �?                      @     �7@     �e@      �?              �?      �?     �F@      �?                       @                       @                       @                33333SK@fffff�@                      �?             �J@      �?       @               @       @       @                       @      �?                fffff�R@ffff��@                                      8@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff&9@     H�@                      �?              <@      �?       @      �?                       @       @       @       @              �?       @333333Z@����̧@      �?              �?      �?     �P@      �?                       @               @       @               @       @              @fffff�P@ffff��@      �?                              $@      �?       @      �?               @                                                       @fffff�S@     �@      �?                              8@              �?               @                               @       @      �?      �?      @�����LI@     #�@                      �?      �?     �Q@      �?       @      �?               @       @               @       @      �?      �?       @     �Z@     �@      �?                              .@      �?       @                                                                      �?       @     �H@     j�@      �?              �?              R@      �?       @      �?               @       @               @       @       @      �?             �Y@33333��@                      �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @     �3@      b@      �?              �?              H@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�����4@     0�@      �?              �?             �Q@      �?       @      �?       @       @       @       @       @       @      �?              �?������\@����� �@                                      @@      �?       @               @                               @       @      �?              @     �R@ffff�ա@                                      =@      �?                       @               @       @                      �?              �?      M@     �@                                      �?      �?              �?                                                              �?       @�����LQ@�����LQ@      �?              �?      �?     �G@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@fffff��@                      �?             �Q@      �?                               @       @       @       @       @       @      �?      �?�����,T@����I�@      �?              �?      �?     �D@      �?       @               @       @       @               @                      �?      �?33333�R@������@                      �?      �?     �Q@      �?       @      �?               @       @       @       @       @       @      �?       @����̌[@�����	�@                      �?              @      �?       @      �?                                       @                      �?       @     �U@     4�@                      �?      �?     �N@      �?       @      �?               @                       @       @              �?       @������X@����z�@      �?                              @      �?       @      �?               @                       @       @              �?       @33333�X@     
�@      �?                              �?      �?              �?                                       @       @              �?       @     PV@     PV@      �?              �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y3@�����mq@      �?                      �?      5@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@     �x@      �?              �?              1@      �?       @      �?               @       @               @       @              �?       @33333�Y@     :�@                      �?      �?      8@              �?               @       @       @               @       @      �?               @������L@     _�@      �?              �?      �?       @      �?       @               @                                                              @�����YL@33333c\@                                      @              �?               @               @                                              @     �A@     �`@      �?                              @              �?               @       @               @                                      @333333E@�����Lb@      �?      �?      �?             �@@      �?       @      �?               @                       @       @              �?        fffff&Y@    ���@                      �?      �?      N@              �?               @               @       @       @       @       @              �?������M@fffff�@      �?                              N@      �?       @      �?               @                       @                      �?        �����yV@3333�J�@                      �?      �?      (@              �?                                       @                      �?              �?     @>@�����w@                      �?              &@      �?       @      �?                                       @       @              �?       @     �W@�����ې@      �?      �?      �?              0@      �?                       @       @                                              �?        fffffFK@�����ȉ@      �?                              <@      �?       @      �?               @                       @       @      �?               @�����Y@ffff� �@                      �?              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�4@fffff�4@                                      .@      �?              �?               @       @               @       @              �?       @     PY@     Ŗ@      �?                              9@      �?       @      �?                                               @              �?       @333333U@������@      �?                              @@      �?       @      �?                                               @              �?        �����iU@�����Ф@              �?                       @      �?       @      �?                                       @                      �?       @33333cU@fffffng@      �?      �?                      E@      �?       @      �?               @                                              �?        fffff�S@33333 �@      �?              �?              8@              �?                               @                                               @�����=@     ��@                                     �M@      �?       @      �?               @       @                                      �?       @     �T@����U�@      �?              �?      �?      D@      �?               @      �?      �?      �?      �?      �?      �?              �?        ffffff4@fffffJ�@      �?              �?      �?     �Q@              �?                       @       @       @       @       @      �?               @�����,N@3333�*�@              �?      �?              �?      �?       @      �?                       @               @       @              �?       @333333Y@333333Y@              �?      �?             �N@      �?       @      �?       @       @       @       @                              �?      �?����̌W@3333s�@      �?      �?                     �Q@      �?       @      �?               @               @       @       @       @      �?       @33333�Z@33333ǽ@                                      8@      �?       @      �?       @                       @                              �?       @fffffU@33333H�@                                      "@      �?               @      �?      �?      �?      �?      �?      �?                             �3@33333�b@      �?                              3@      �?              �?               @       @                                      �?       @     �S@�����K�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �3@33333`@      �?              �?              E@      �?       @               @                                              �?              �?�����L@3333���@      �?                             �A@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @3333334@33333c�@      �?                             �@@              �?                       @                       @              �?      �?       @����̌C@     t�@      �?              �?      �?      <@      �?              �?                       @               @                               @�����\U@������@      �?              �?              1@              �?               @               @                                              @333333A@     ��@                                      F@              �?                               @               @       @      �?      �?       @fffff�H@     ��@                              �?      5@      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@33333C|@      �?      �?      �?             �Q@      �?       @               @       @       @       @       @       @       @      �?      �?33333#V@    ���@                                      $@      �?              �?       @                               @                      �?      @�����,U@fffff �@              �?                      G@      �?       @                               @       @               @      �?      �?      �?fffffFQ@3333�n�@                                      >@      �?       @                       @       @               @              �?      �?      �?�����<Q@�����ڟ@                              �?      :@              �?               @                       @               @                      @fffff�F@     �@                                      <@      �?       @                                       @                              �?      �?33333sK@�������@                      �?      �?     �M@      �?       @               @               @       @       @               @      �?      @�����S@    ���@                                      .@      �?       @                                                                      �?      @ffffffH@����̀�@      �?                             �B@      �?              �?                                                              �?      @fffff�Q@������@      �?      �?                      P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����4@33333��@      �?              �?      �?       @      �?                                                                                        33333SF@fffffw@      �?                      �?      @      �?       @      �?               @                       @       @              �?       @�����lY@������v@      �?                              �?      �?                                                                                       @fffff�F@fffff�F@                                       @      �?                       @       @               @                      �?                �����M@     T}@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @����̌3@33333`@                      �?              L@      �?              �?       @               @                               @                33333T@ffff���@      �?                               @      �?              �?       @       @                       @       @                       @�����Y@     �h@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����L3@�����L3@      �?      �?                      $@      �?       @      �?                                       @       @              �?       @fffff�W@������@                                     �E@      �?              �?               @       @               @                      �?       @������V@33333�@              �?      �?              O@      �?                       @               @       @       @       @       @      �?      �?������S@    �Ӳ@                      �?               @      �?              �?               @       @               @       @                       @�����IY@33333W�@      �?      �?                     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����L4@333331�@                              �?      �?      �?              �?       @                                                      �?      @ffffffR@ffffffR@                                      B@      �?                       @       @       @       @       @              �?      �?      @fffffS@3333�\�@      �?              �?      �?      �?      �?              �?                                                              �?       @      Q@      Q@                                      @      �?              �?                                                              �?      @     PQ@fffff&z@      �?      �?      �?             �D@      �?       @      �?       @               @                                      �?             �T@������@      �?              �?      �?      ?@              �?               @                       @                                        33333�A@     ֐@                      �?              5@              �?               @                                                               @     �<@����̪�@      �?              �?      �?     �H@              �?               @                                       @              �?       @������C@�������@      �?                      �?      �?      �?       @      �?                       @               @       @              �?       @     �X@     �X@      �?              �?              B@      �?               @      �?      �?      �?      �?      �?      �?      �?              @      4@     ք@      �?              �?      �?     @Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?              :@33333�@      �?                              &@      �?              �?       @               @                                      �?             �S@33333݈@              �?                      @      �?       @      �?                                                              �?       @����̜R@33333gr@      �?                              "@      �?              �?                                                              �?       @     �Q@33333��@                      �?             �G@      �?                       @               @               @              �?      �?      �?33333�P@ffff暧@              �?                      @      �?                       @       @               @                                      �?33333�M@������q@                                      @      �?              �?       @       @       @       @               @              �?        ������X@�������@                      �?      �?     �B@      �?       @      �?               @       @                       @              �?       @������W@3333���@                      �?      �?      Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        �����Y3@�����2�@      �?      �?      �?      �?      P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        ffffff8@�����2�@      �?                              �?      �?              �?                                                              �?       @ffffffQ@ffffffQ@      �?              �?      �?      L@              �?               @       @               @       @              �?      �?      @      J@����̉�@              �?      �?             �G@      �?       @               @       @       @                                      �?      �?������P@     h�@                                      R@      �?       @      �?               @       @       @       @       @       @      �?        fffff�[@    �L�@              �?                      2@      �?              �?                       @                       @              �?       @�����<U@�������@                      �?              :@      �?       @      �?               @                                                        33333�S@33333�@                                      .@              �?               @       @       @       @                      �?              @33333�F@�������@                      �?      �?      0@      �?       @      �?               @                                              �?      �?������S@�����ϓ@                                      (@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@fffffNp@                      �?              R@      �?       @      �?               @       @       @       @       @      �?              �?�����I[@�����m�@                                      �?      �?                                                                              �?       @fffff�F@fffff�F@      �?                              R@      �?       @      �?       @       @       @       @       @       @       @                �����Y\@�����@                      �?              G@              �?                                               @       @              �?       @������E@fffff_�@      �?                              �?      �?                               @                                              �?       @     `I@     `I@              �?                      �?      �?       @      �?                                                              �?       @fffffR@fffffR@      �?              �?              Q@      �?              �?               @               @       @       @      �?      �?       @33333Y@����Yb�@      �?              �?             �P@      �?       @      �?               @               @       @       @      �?      �?       @33333Z@     �@      �?                      �?      C@      �?       @      �?               @                                              �?      @fffffvT@fffff��@      �?      �?      �?              R@      �?       @               @       @       @               @       @       @      �?      �?fffffU@ffff�]�@      �?                             �@@      �?       @      �?       @                                              �?                fffffT@�����V�@      �?      �?                      3@      �?       @      �?               @                       @                      �?       @�����V@33333��@              �?                      .@      �?              �?                                       @       @              �?       @     �V@33333�@      �?                             �C@              �?                               @       @                      �?              @fffff�A@�����t�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff&4@fffff&4@      �?              �?      �?     �B@      �?                       @               @       @                      �?      �?      @     `M@333336�@                      �?             �Q@              �?               @       @       @       @       @       @       @                33333#P@ffff昱@      �?              �?      �?      P@      �?       @      �?                       @                       @      �?              �?     �V@ffff&��@      �?      �?                      �?      �?              �?                                                              �?       @     pQ@     pQ@      �?                             �O@      �?       @      �?               @               @       @       @                       @�����YZ@333339�@                                      (@      �?       @      �?                                       @       @              �?       @����̌W@fffffX�@                      �?      �?      (@      �?               @      �?      �?      �?      �?      �?      �?                        ffffff3@33333�h@              �?                     �H@      �?       @      �?                       @                       @              �?      �?fffff�V@����٣�@              �?      �?              @              �?                       @                                              �?       @     �>@fffff�T@                      �?             �L@      �?       @      �?       @                               @       @              �?       @������X@����y�@                      �?      �?      @              �?               @                                                              �?33333�=@������V@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�2@������[@                      �?              R@      �?       @               @       @       @       @       @       @       @      �?       @�����W@������@              �?                     �F@      �?              �?       @       @               @                              �?        �����lU@33333��@                                      �?      �?       @      �?                                               @                      @33333sU@33333sU@                                       @              �?                       @                       @       @                       @33333�I@333333X@                      �?      �?      7@      �?                       @       @       @       @                      �?      �?      @     �P@33333��@      �?              �?              Q@      �?       @               @       @       @       @       @       @       @      �?      �?33333�V@����ٞ�@      �?              �?              C@      �?              �?       @       @                                              �?       @������S@������@      �?      �?      �?             @Q@              �?                               @                              �?      �?      �?������=@�������@                      �?      �?     �B@      �?               @      �?      �?      �?      �?      �?      �?                       @�����Y3@     ^�@      �?      �?                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����4@      �?                             �O@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �4@�������@                                     �K@      �?       @      �?       @               @                              �?      �?      �?     U@������@                      �?             �L@      �?       @      �?               @       @       @       @       @      �?      �?        �����Y[@3333�l�@                                      *@      �?       @      �?                                               @              �?       @�����|U@�������@              �?      �?             �Q@      �?              �?               @       @                       @       @              �?�����\V@    @#�@      �?              �?             �P@      �?       @               @       @       @       @                       @              �?������Q@����E�@      �?              �?             @Q@      �?       @      �?               @               @       @               @      �?      @�����W@���̌<�@      �?                              @      �?       @                                       @               @                      @33333cP@fffff�m@      �?                              �?      �?                                       @       @       @       @              �?       @     �R@     �R@                                      $@      �?                                       @       @                                       @      K@     8�@      �?                             �@@      �?                               @       @               @                      �?      �?������P@����̊�@                      �?      �?      L@      �?              �?                                       @       @      �?                �����9V@     h�@      �?              �?      �?     �@@      �?                               @       @       @       @       @       @              �?fffff�T@33333V�@      �?                              (@      �?                               @                                              �?        fffff�H@fffff��@      �?              �?      �?      &@      �?                                       @               @                      �?        33333�M@     Z�@                      �?             �B@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ������3@     l�@      �?      �?      �?      �?      Q@      �?               @      �?      �?      �?      �?      �?      �?      �?                     �3@33333��@                                      >@      �?               @      �?      �?      �?      �?      �?      �?       @              �?ffffff3@     �@      �?              �?      �?      (@              �?                       @               @                                      @     �A@     {@      �?              �?      �?      L@      �?       @      �?       @       @       @       @       @       @       @              @fffff�\@ffff槹@      �?                              @      �?                                       @       @                                       @33333L@333337r@                                      .@      �?               @      �?      �?      �?      �?      �?      �?                             �3@����̔r@                                      .@      �?              �?       @                               @                               @����̌U@�����ؓ@      �?              �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff&9@�������@      �?              �?      �?     �M@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@     ��@      �?                      �?      ;@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?������9@fffff��@                      �?              �?      �?              �?                                       @                      �?        fffff�S@fffff�S@      �?              �?      �?      C@      �?                       @               @       @       @       @       @              �?     @T@������@              �?      �?             �C@      �?              �?       @       @                       @       @      �?              @fffff�X@ffff�K�@                                      9@      �?                       @       @       @       @       @              �?              @33333�R@33333�@      �?      �?                      0@              �?                       @                       @                      �?      @     �C@�����>�@                                      &@      �?                                                                              �?      @33333SF@     �}@                                      (@              �?               @               @       @               @       @              @������H@�����@�@      �?                              &@      �?              �?               @                                                       @����̼R@     |�@                      �?              �?      �?              �?                                       @                               @33333�S@33333�S@      �?      �?                      ,@      �?       @      �?                                                              �?       @����̼R@     3�@      �?              �?      �?     �J@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?3333334@�������@      �?      �?      �?              @      �?              �?                       @               @       @              �?       @     �W@     �@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?�����]@    ���@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?             @:@33333�@      �?              �?      �?      @      �?              �?                                                              �?       @33333sQ@������w@      �?      �?                     @P@      �?       @      �?       @               @       @       @       @       @      �?       @fffff�[@ffff&N�@      �?      �?                      �?      �?                                                                                       @����̌F@����̌F@      �?                              D@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @������8@�����o�@                      �?      �?       @      �?              �?                                                              �?       @������Q@     �`@                              �?       @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@�����\e@                      �?      �?     �C@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ������3@fffff��@                              �?      @              �?               @                                                              @������=@fffff>i@      �?                              �?              �?                                                       @                       @33333�A@33333�A@              �?                      �?      �?              �?                                                              �?       @     PQ@     PQ@                      �?      �?      J@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����9@     ٓ@      �?      �?      �?              $@      �?              �?               @       @       @       @                      �?      @      W@�����0�@      �?                              (@      �?       @      �?                                       @       @                       @33333�W@33333V�@                      �?              4@      �?              �?                                                              �?        33333sQ@fffff�@      �?              �?      �?      9@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     �9@����̴�@                      �?      �?     �Q@              �?               @       @               @       @       @       @                ������M@ffff��@                              �?      �?              �?                                                                              @33333�8@33333�8@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                       @     �3@     �3@      �?                             �M@      �?       @                               @                               @              �?33333K@����LX�@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                        33333�3@33333�3@      �?                              P@      �?       @               @       @       @       @       @              �?               @     PT@���̌��@                                      6@      �?              �?               @                               @              �?      @33333U@�������@      �?              �?              G@      �?                       @       @       @       @                       @              @�����iP@����LΧ@      �?      �?      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?33333s9@�������@      �?              �?      �?      <@      �?       @                       @                               @                       @�����P@�����(�@                                      E@      �?                                       @       @               @       @              �?     �P@    ���@                                     �J@              �?               @       @       @       @       @              �?      �?       @������J@fffff~�@      �?      �?      �?              =@      �?       @      �?                       @               @       @              �?       @     �X@����Lx�@                      �?      �?     �E@      �?                                                       @                               @33333L@�������@      �?      �?                      1@      �?              �?               @       @               @       @              �?       @33333sY@�����a�@      �?      �?      �?              =@      �?       @      �?                                       @       @              �?       @����̜W@����L��@      �?                      �?      3@      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?�����8@33333s{@      �?      �?                      @      �?       @      �?                                                                      @     pR@33333	�@              �?      �?             �G@      �?       @      �?                       @               @       @                       @������X@33333��@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@�����)S@                      �?              P@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333s3@�����&�@      �?                              F@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����4@     j�@      �?      �?                     �F@      �?                       @               @                       @      �?              �?�����YO@     ϥ@      �?                              (@              �?               @       @               @       @                      �?        �����yI@     �@      �?              �?              ?@      �?       @      �?               @       @               @                               @33333sW@     ��@                                     �C@              �?                       @       @       @                                        ����̌D@33333��@                                      =@      �?               @      �?      �?      �?      �?      �?      �?                      �?�����Y3@�����̂@                                      <@              �?                               @                                      �?      @     �=@�������@                      �?      �?      5@      �?              �?               @                                              �?        33333�R@�����v�@              �?      �?              6@      �?       @               @       @               @                              �?      @fffff�O@33333��@                      �?      �?     �A@              �?               @                       @       @               @      �?      �?�����,G@33333��@      �?              �?      �?     �O@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@fffff�@      �?                              �?      �?                                               @                                      �?     �H@     �H@      �?              �?      �?     �E@      �?       @      �?       @               @       @                      �?      �?      �?     �V@�����[�@      �?                             �H@      �?       @                                       @       @               @      �?        ������P@     ��@      �?                              ;@      �?              �?                                                              �?      @33333CQ@     �@                                      ,@      �?              �?                                       @       @              �?      @33333sV@fffff��@                                      @      �?              �?               @                       @       @      �?      �?      @33333�W@�����˃@                                      N@      �?              �?               @       @               @       @       @      �?       @������X@����5�@      �?              �?      �?      P@              �?               @               @       @       @       @       @      �?        fffffN@ffff�
�@      �?                              �?      �?              �?                                       @                      �?       @33333�S@33333�S@      �?                              @@      �?              �?                               @       @       @              �?       @�����X@�����ި@                      �?      �?      7@      �?               @      �?      �?      �?      �?      �?      �?       @                ffffff4@     �}@                                      C@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����L4@fffff8�@                                     �A@      �?                       @       @       @                                               @fffffFN@fffff��@                      �?      �?     �Q@      �?       @               @       @       @       @       @       @       @              @33333�V@    ���@                      �?      �?      8@              �?               @       @       @       @               @       @      �?      @     @J@�������@      �?              �?      �?      2@      �?                                       @                       @                       @������L@�������@      �?      �?      �?               @      �?       @      �?                                       @                      �?      @fffff�U@33333�c@      �?              �?      �?      E@      �?                       @       @                                                      @     @K@����L��@      �?                              C@      �?       @      �?               @       @                       @              �?      �?fffff�W@fffff֬@      �?              �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�3@�����2�@      �?                              @      �?                                                                                      @������F@fffff�a@                                      �?      �?       @      �?               @                                              �?      @�����T@�����T@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?                      @������3@�����Yf@                                      �?              �?                                               @                      �?       @�����YA@�����YA@      �?                              "@              �?               @       @       @                              �?              @fffff�C@     Pw@      �?                              4@      �?       @      �?                               @       @       @              �?      @33333�X@����̿�@      �?      �?                      5@      �?              �?                       @               @       @              �?        333333X@33333��@              �?      �?              6@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                ������9@fffff&�@      �?              �?      �?      9@      �?                       @                       @                                       @fffff&K@33333C�@                      �?              @      �?                       @                                                      �?        fffff&I@�����1v@                      �?             �C@              �?               @               @               @       @                       @33333�K@3333��@      �?              �?              @              �?                                                                      �?       @33333�8@�����Y@              �?      �?             @P@      �?       @      �?               @       @               @       @      �?      �?       @     �Z@�����C�@      �?                              4@      �?              �?       @       @       @       @       @       @              �?        �����[@fffff7�@      �?              �?      �?      1@      �?              �?                                       @                               @fffff6T@fffff�@      �?              �?              1@      �?                       @       @                               @      �?              @333333P@fffff^�@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @ffffff4@ffffff4@      �?                              4@      �?                               @                                              �?      @fffff�I@�������@                      �?             �B@              �?               @                       @       @               @               @33333�F@fffff�@      �?              �?             �N@      �?       @                       @       @               @       @       @                �����9T@    �D�@      �?                      �?     �C@              �?                               @       @       @       @      �?                �����lK@fffff�@                                     �P@      �?                       @       @               @                      �?              �?     @N@     <�@              �?      �?             �A@      �?       @      �?                       @               @       @                        33333�Y@������@                                      P@      �?       @               @       @       @       @       @       @       @      �?      �?������U@����B�@      �?              �?      �?      3@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@     �u@                                      �?      �?       @      �?                                       @       @              �?       @fffffvW@fffffvW@                      �?      �?       @      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@�����Dd@                      �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @3333333@������@                                      &@      �?       @      �?                       @               @       @              �?       @     0Y@     ��@              �?                      :@      �?              �?                                       @       @              �?       @     �V@�����_�@                      �?              �?      �?                                                       @                              @������K@������K@                                      @      �?               @      �?      �?      �?      �?      �?      �?       @              @����̌3@�����_@              �?      �?             �Q@      �?       @      �?       @                                               @      �?      �?�����,T@     ,�@      �?                             �A@      �?                       @       @       @                              �?              @������N@����̔�@      �?              �?      �?      7@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@fffff�z@      �?              �?             �F@      �?       @      �?       @               @                                      �?      @33333#U@ffff��@                      �?               @      �?               @      �?      �?      �?      �?      �?      �?                        ������3@      J@      �?              �?             �O@      �?               @      �?      �?      �?      �?      �?      �?       @              @     @3@�����V�@                                      B@      �?       @                       @               @               @      �?      �?      @����̬Q@ffff柣@                                      @      �?              �?                                                              �?       @������Q@������p@      �?              �?      �?      R@              �?               @               @       @       @               @              @33333sH@     ��@      �?              �?             �Q@              �?                       @                       @       @       @               @����̬H@    �v�@      �?              �?             �Q@      �?       @      �?       @       @       @       @       @       @       @              �?33333�\@ffff&�@      �?                             �P@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @33333s3@����̯�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?              �?        33333�3@�����e@      �?                             �F@      �?       @      �?               @                       @       @              �?      �?fffff6Y@     ��@                      �?      �?      M@              �?               @               @       @       @       @       @              @     �M@3333�P�@      �?      �?      �?              @@      �?              �?                                               @              �?      �?33333T@����f�@                      �?      �?     �B@      �?                       @       @                       @       @      �?                fffff�R@�����Ť@      �?              �?              R@      �?       @                       @       @               @       @       @                ������T@����L��@              �?                      ,@      �?       @      �?                                                              �?       @33333�R@     !�@      �?                      �?      :@              �?                       @                       @              �?      �?        ������C@     ��@      �?              �?              "@      �?       @      �?       @                                       @              �?       @33333V@fffff
�@              �?                     �O@      �?       @      �?                       @                       @              �?        ffffffV@����̢�@                                      $@              �?               @       @       @                                                �����YD@�����|@                      �?      �?     @Q@      �?       @      �?       @       @       @       @       @       @       @              �?     P\@ffff&׾@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @3333333@33333�c@      �?                              "@      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@     Pf@                              �?      .@      �?              �?               @                               @              �?        �����yU@33333֓@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @������3@33333�]@                                       @      �?       @      �?                                               @              �?       @�����lU@�����9e@                                      =@      �?       @      �?                                                              �?       @����̌R@     %�@      �?      �?                      N@      �?       @               @       @                               @      �?      �?       @     �Q@���̌�@                                     �D@      �?               @      �?      �?      �?      �?      �?      �?                       @33333s4@�����<�@      �?      �?      �?              @      �?       @      �?               @       @               @       @              �?       @�����yZ@fffff�t@      �?                             �@@      �?       @                       @                                              �?        33333SK@������@                                      @      �?       @                                                                      �?      @33333SI@������b@                      �?      �?     �I@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�3@     �@      �?                              �?      �?              �?                                                              �?       @�����yQ@�����yQ@      �?                              $@      �?              �?                                       @       @              �?       @     `V@�������@              �?                      �?      �?              �?                                                              �?       @������Q@������Q@      �?              �?      �?      @      �?              �?                                                              �?        �����|Q@     ��@      �?              �?              D@      �?       @      �?               @                       @       @              �?       @33333SY@�����@      �?                              �?      �?       @      �?                                                              �?       @������R@������R@              �?                      J@      �?       @               @               @                               @                ������M@    �>�@              �?                      �?      �?              �?                                                              �?       @ffffffQ@ffffffQ@      �?              �?      �?     @P@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@fffff2�@                                       @      �?       @      �?                                       @       @              �?       @      X@������e@      �?              �?             �P@      �?       @                                       @               @                       @������O@�������@                      �?               @      �?              �?                                                              �?       @fffff�Q@     ^@      �?              �?      �?      3@              �?               @       @                                              �?      @�����yA@������@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @����̌3@����̌3@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @      3@������S@                      �?              >@      �?               @      �?      �?      �?      �?      �?      �?                        fffff�3@�����~�@      �?              �?      �?     �Q@      �?       @               @       @               @                      �?      �?      �?fffff�P@3333���@                              �?      ?@      �?       @      �?                                       @                      �?      �?33333�U@������@      �?      �?      �?              H@      �?       @      �?                       @                       @              �?      �?33333�V@    ��@      �?                              3@              �?                                                                      �?        fffff&9@�����E}@                                      $@      �?               @      �?      �?      �?      �?      �?      �?              �?       @3333335@������k@              �?      �?              R@      �?       @      �?               @       @               @       @      �?              �?     @Z@������@      �?                             �A@      �?       @      �?       @       @       @       @                              �?      @     0X@����̖�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?      �?              @3333335@fffffJ@      �?              �?              H@      �?       @                       @       @                       @      �?      �?      �?33333�Q@     ��@      �?      �?      �?              ;@      �?              �?                                                              �?       @33333�Q@�����_�@      �?                              2@      �?                       @               @       @       @                      �?       @fffffQ@33333O�@                                       @      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff3@fffff�N@      �?                              &@      �?                                       @               @       @              �?       @fffffVQ@     B�@      �?                             @Q@      �?       @      �?       @       @       @               @       @       @      �?      �?33333�[@    ��@      �?      �?                      8@      �?              �?                                                                      �?     �Q@fffff�@                              �?      5@      �?                       @               @                       @      �?              @fffff6P@33333�@      �?                              &@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?33333s4@������m@                                      @      �?                       @                                                      �?        fffffFI@�����tm@                      �?      �?     �K@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?fffff�9@     ��@                      �?      �?      (@      �?               @      �?      �?      �?      �?      �?      �?       @                �����L4@     l@      �?              �?      �?      A@      �?       @      �?                       @                       @              �?      �?33333�V@     2�@      �?                              �?      �?                                       @                                      �?      @33333�H@33333�H@      �?      �?                       @      �?       @      �?                       @               @       @              �?       @fffff&Y@33333��@      �?              �?      �?      R@      �?       @               @       @       @       @                       @              �?fffffR@ffff���@                      �?      �?      R@      �?       @                       @               @       @       @       @      �?       @����̼S@ffff&b�@                                     �O@      �?                                       @                       @      �?              �?fffffFM@     _�@                                      �?      �?                                                                                      �?������E@������E@              �?                      @      �?       @      �?               @                                              �?       @������S@������i@      �?              �?      �?      .@      �?              �?       @                                                              @fffff�R@33333��@                      �?      �?      1@      �?              �?       @                       @       @                               @fffff�V@����̙�@                                      @      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @fffff�7@     `X@      �?              �?              @              �?                                       @                              �?       @fffff�=@     W@      �?              �?               @      �?                               @               @               @              �?      @�����P@������a@      �?      �?      �?              Q@              �?               @       @       @                               @      �?       @������D@    �+�@      �?                             �L@      �?       @      �?                               @       @               @      �?      �?����̜V@�����m�@                      �?              ;@      �?       @      �?                       @                       @                        ������V@������@      �?      �?      �?             �J@      �?       @      �?               @       @               @       @              �?       @fffff�Y@    �m�@                      �?               @      �?              �?                                                              �?       @����̬Q@fffff�a@                      �?             �Q@      �?       @               @               @       @                       @              �?33333SP@    ���@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�4@     0\@      �?      �?                      4@      �?                       @                       @                      �?              @      K@������@      �?              �?      �?      C@      �?       @      �?                       @       @       @               @      �?        ������W@    �@�@      �?              �?      �?      D@      �?              �?                       @               @              �?      �?       @33333CU@����L7�@                                     �E@      �?       @      �?       @       @       @       @       @       @       @              �?33333�\@�����@      �?      �?      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333�7@�����p�@      �?      �?      �?             �P@      �?       @      �?                                       @       @              �?      �?������W@     ��@      �?              �?              <@      �?                       @       @               @                                      @33333sN@������@                      �?      �?      8@      �?       @               @       @                       @       @      �?               @������S@�������@                      �?              L@      �?       @      �?       @       @       @               @       @      �?                33333s[@ffff�ݷ@      �?              �?             �P@      �?              �?       @       @                               @      �?      �?      �?fffff�V@ffff&��@                                      @      �?              �?                       @       @                                      �?fffffT@�����1k@      �?              �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                fffff&9@fffffS�@                      �?      �?      H@      �?       @                       @               @       @       @       @               @������S@�����<�@      �?                               @              �?                                                                      �?       @�����9@�����,L@      �?              �?      �?      ?@      �?       @                                                       @                        ������M@     ��@      �?                              J@      �?                       @       @                       @               @      �?      �?     �O@ffff��@                      �?      �?     �P@              �?                       @       @       @       @       @       @      �?       @fffff�M@ffff��@                                      D@      �?       @                               @       @       @       @      �?      �?      @     0T@����L�@                      �?             �M@      �?               @      �?      �?      �?      �?      �?      �?       @                ffffff2@fffff��@      �?                              @      �?              �?                                                              �?      @33333�Q@����̌k@                                      7@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              �?������8@�����:�@              �?      �?              ;@      �?       @                       @       @       @       @       @                       @fffff�T@fffff�@      �?      �?      �?              0@      �?       @      �?                       @               @       @              �?       @     �X@33333Θ@      �?                      �?      �?              �?                                                                              @3333338@3333338@                      �?      �?      2@      �?                                       @       @                      �?      �?      �?333333K@������@      �?                              @      �?       @      �?                                                                      @     �R@33333#j@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?      �?fffff�\@fffff��@      �?              �?              6@      �?              �?                       @               @       @              �?      �?����̬W@������@      �?                              1@      �?                       @       @                                              �?      �?     �K@333331�@                                      @      �?                                               @                              �?        33333�H@������p@      �?              �?      �?      @@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333�2@�����/�@                                      D@      �?       @      �?                       @       @       @       @      �?      �?      �?�����|Z@33333�@                      �?      �?      ?@      �?       @      �?               @                               @              �?       @������V@ffff�f�@                                     �J@      �?              �?       @       @       @       @               @       @              @     �X@    @0�@      �?      �?      �?             @Q@      �?       @      �?       @               @       @       @       @      �?      �?      @33333�[@������@      �?      �?                      J@              �?                       @                       @       @              �?       @33333�H@������@                      �?      �?      B@      �?                       @                                                              �?fffff�I@     \�@                                      B@      �?                       @       @       @       @       @       @      �?                fffffvU@����w�@      �?              �?              "@              �?                                                              �?                �����8@�����<p@                                      "@              �?                       @                               @                       @     `D@fffffvv@                      �?             @Q@      �?       @      �?                       @       @       @       @       @                fffffVZ@ffff�H�@                                     �D@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @     �3@�����7�@                                      "@      �?              �?                                       @       @              �?      @�����V@����̤�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                       @fffff�4@fffff�4@              �?                      &@      �?       @               @                                                      �?       @������K@fffff&�@      �?              �?             �P@      �?       @      �?               @                       @              �?      �?        �����V@����L��@              �?      �?             @Q@      �?              �?       @       @                               @      �?              �?33333�U@���̌��@                      �?             �Q@      �?       @      �?                                       @       @       @      �?        �����lW@����Y��@      �?              �?      �?      A@      �?              �?                                       @                               @33333�S@������@      �?                      �?     �J@      �?                       @       @               @                      �?              �?�����lO@     ��@      �?              �?               @      �?       @      �?                                               @              �?        �����iU@�������@              �?                      "@      �?       @      �?                                                              �?       @33333�R@33333w�@                      �?              O@      �?              �?       @               @       @       @       @      �?      �?       @33333Z@ffff�չ@              �?                      P@      �?       @      �?       @               @       @       @       @              �?        �����<[@����Lǻ@              �?                      K@      �?       @      �?               @                                              �?       @     �S@    @�@                      �?      �?     �L@      �?       @               @               @       @       @       @       @      �?       @      U@fffff�@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?              �?      �?������4@     �t@      �?                               @      �?              �?               @                                              �?       @     �R@�����b@                                      @              �?                                                                                �����9@fffff�g@                      �?      �?     �G@              �?               @       @       @               @       @       @      �?      �?      N@����L��@                      �?             �G@      �?       @       @      �?      �?      �?      �?      �?      �?      �?               @fffff�:@fffff��@                                      =@      �?              �?                                       @                      �?       @������S@����L��@                                      2@      �?       @      �?                               @               @              �?       @fffff�V@     3�@      �?                      �?      =@              �?               @       @       @       @                              �?      @     �F@�����i�@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @              �?�����lV@����Lø@                                      �?      �?              �?                               @       @       @              �?       @fffff�W@fffff�W@      �?                              R@      �?               @      �?      �?      �?      �?      �?      �?       @                ������3@fffffh�@                                      @              �?                                                                      �?       @33333s8@fffff�U@      �?      �?                     �H@      �?       @      �?                                       @       @              �?       @�����X@    @n�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                        fffff&4@     P`@      �?                             �B@      �?       @      �?                               @       @       @                        33333�X@����'�@      �?      �?                     �P@      �?       @               @       @               @                       @      �?        33333#P@������@                                      I@      �?       @      �?       @       @               @       @       @       @      �?       @�����i[@ffff&��@      �?      �?      �?              P@      �?       @      �?                       @       @       @       @       @               @fffff�Y@3333s��@      �?                              @      �?              �?                       @                                              @������R@fffff�@      �?                              G@      �?               @      �?      �?      �?      �?      �?      �?       @              �?3333333@33333a�@                      �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@33333SN@      �?              �?      �?      N@      �?       @      �?               @               @       @       @              �?             �Y@3333�Q�@                      �?      �?     �F@              �?               @                               @       @              �?        33333sI@3333�;�@      �?              �?      �?      8@      �?       @               @               @       @       @       @      �?      �?      @333333U@     �@      �?                              @      �?       @      �?                       @               @                      �?      �?fffffVV@����̾�@                      �?              Q@      �?       @               @                       @                      �?                      M@fffff�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@     @4@              �?      �?              @      �?       @      �?       @                               @       @              �?       @fffff�X@fffff�u@                                      I@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @�����Y3@     $�@                      �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?        ����̌\@ffff�+�@              �?                      �?      �?       @                                                                              @fffffFI@fffffFI@      �?                              G@              �?               @                                              �?      �?             �>@33333E�@                                      �?      �?              �?       @                               @       @              �?       @fffff�W@fffff�W@      �?      �?      �?              *@      �?              �?               @               @               @              �?        33333CV@fffffE�@                              �?     �Q@      �?       @               @       @               @                       @               @     �P@    ��@                                       @      �?       @               @       @       @                                      �?             `P@33333�@      �?              �?             �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������9@������@      �?                             �L@              �?                               @       @       @       @       @              �?����̬J@����$�@      �?              �?      �?      @      �?                                       @                                      �?       @33333I@�����e@                                      @      �?       @      �?               @                                              �?      @33333T@33333Ct@                                      �?      �?              �?                                                                        �����lQ@�����lQ@      �?      �?      �?              I@      �?       @      �?       @               @               @       @       @      �?      �?33333CZ@����L+�@                                      1@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff&4@fffffv@      �?              �?              @      �?       @                               @               @                               @ffffffP@33333Co@      �?                      �?      A@      �?       @      �?       @       @                       @       @      �?      �?       @33333�Y@������@      �?              �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?              �?       @      4@����� r@              �?                      O@      �?       @      �?                                       @              �?               @�����U@ffff&_�@              �?      �?             �L@      �?       @      �?               @       @                       @                      �?     �W@3333�>�@      �?              �?               @      �?       @      �?                       @               @                      �?       @������V@fffffne@                                      $@      �?       @      �?       @                               @       @              �?       @����̬X@     j�@      �?                              B@      �?                       @               @       @       @       @              �?      �?������S@ffff�M�@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@fffffFU@      �?      �?      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                ������8@     ��@      �?      �?      �?             �I@      �?       @      �?       @               @                       @      �?      �?        �����iW@ffff&�@                                      G@      �?              �?       @       @       @               @              �?      �?      �?������W@333338�@      �?              �?      �?      R@              �?               @       @       @       @       @       @       @      �?        �����iP@    �8�@                      �?              :@      �?              �?                               @               @                      �?�����yU@ffff�(�@              �?                       @      �?              �?               @                       @                      �?        33333�T@fffffvd@      �?              �?              6@      �?                       @                       @                      �?      �?      �?      L@�����0�@      �?                              B@      �?       @      �?                                               @              �?       @     0U@����Lԧ@              �?                     �L@              �?                       @       @               @       @              �?       @     �K@����,�@                      �?              L@      �?       @      �?               @       @       @                                       @33333�V@�������@                      �?               @      �?       @      �?                                               @              �?       @�����9U@������@                      �?              D@      �?       @      �?                               @                              �?      �?fffff�S@3333�m�@              �?      �?      �?      L@      �?                       @                       @       @       @       @      �?      �?fffff&R@3333��@              �?                      *@      �?                               @       @                                      �?       @ffffffK@fffffچ@                      �?              �?      �?              �?                                                              �?       @�����<Q@�����<Q@                                       @      �?              �?                                       @                      �?              T@����̄�@      �?      �?      �?              6@      �?              �?                                       @       @              �?             pV@�����K�@      �?      �?                      @      �?              �?                                       @                      �?       @������S@fffffNp@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@�����Y4@                              �?      2@              �?                                                       @              �?       @     �A@     H�@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @3333333@3333333@                      �?      �?      @@      �?                       @       @       @       @               @       @              @ffffffR@3333��@      �?      �?      �?             �D@      �?       @      �?                       @               @       @              �?       @33333�X@����L��@              �?      �?             �Q@      �?       @      �?               @               @       @       @      �?      �?        33333cZ@����Y�@      �?                              @      �?                                       @               @       @              �?       @33333�Q@fffff�u@      �?                             �C@              �?                                       @               @              �?       @�����LD@     Z�@      �?              �?      �?      <@      �?       @      �?                                       @       @      �?                �����W@����L�@                      �?      �?      =@      �?              �?                                       @       @              �?      �?33333�U@    �{�@                      �?              @      �?       @      �?               @                               @              �?      �?     �V@fffff^n@                                      .@      �?               @      �?      �?      �?      �?      �?      �?                        ffffff3@�����r@                                     �I@      �?              �?                                       @       @      �?              �?33333�U@ffff�{�@                                       @      �?                       @                                                      �?       @������H@������v@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����4@      �?              �?      �?     �H@              �?                       @                       @       @      �?      �?        fffff�I@    �ڣ@                                       @      �?       @               @                       @               @                       @������Q@33333��@              �?                      ?@      �?       @      �?               @                       @       @              �?       @������X@����L�@      �?              �?             �Q@      �?       @      �?               @       @       @               @       @      �?        ����̬X@ffff�ʺ@                      �?      �?      �?      �?              �?                                       @                      �?      @33333T@33333T@      �?                              1@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff&3@33333wu@      �?              �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@33333g�@      �?                      �?      =@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@fffff��@                      �?              :@      �?                               @       @       @       @       @                        �����yT@����=�@                      �?      �?      J@      �?       @      �?                       @               @       @      �?                     PY@������@      �?              �?      �?      C@      �?               @      �?      �?      �?      �?      �?      �?                       @������3@fffffj�@      �?              �?             �P@      �?       @      �?               @       @                       @       @      �?       @�����IW@33333�@                      �?      �?      >@      �?                               @       @       @       @       @       @                333333T@�������@              �?                      :@      �?       @      �?       @       @                               @              �?       @     �W@fffff��@                      �?      �?      >@      �?               @      �?      �?      �?      �?      �?      �?      �?                ����̌3@     �@                                      A@      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@�����	�@      �?                              8@      �?              �?               @       @                       @              �?       @33333cV@����L�@      �?              �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?������3@������@      �?      �?      �?             �P@      �?       @      �?                               @       @       @              �?      �?33333Y@ffff�׺@                                      2@      �?              �?       @                                                      �?       @������R@�������@                      �?      �?      J@      �?       @      �?               @       @               @              �?      �?      �?������W@ffff&p�@                      �?      �?      H@      �?               @      �?      �?      �?      �?      �?      �?       @              @����̌3@����̚�@      �?      �?      �?              R@              �?               @       @       @       @       @       @       @      �?        ����̌O@���̌M�@      �?                              4@      �?       @                       @               @       @              �?      �?       @�����,Q@����� �@      �?              �?             �G@      �?       @      �?               @                                      �?      �?       @������S@3333���@      �?      �?                      Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?      4@     Е@      �?                             �I@      �?       @      �?               @                                                             @T@    ��@                              �?      6@      �?               @      �?      �?      �?      �?      �?      �?              �?       @����̌4@�����]}@      �?              �?      �?      G@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        3333334@�����l�@      �?                               @      �?                                                               @              �?      �?     `K@�����`{@                                     �G@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff&4@�����X�@      �?      �?                      �?      �?              �?                                                              �?       @������Q@������Q@                                      E@      �?              �?               @       @       @       @       @              �?        33333�Y@    ��@              �?      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff�\@�����>�@      �?                              :@      �?       @      �?       @       @                       @                      �?      �?�����W@�����[�@                      �?             �O@      �?       @      �?               @       @       @       @       @       @      �?             P[@fffff��@                                      @      �?              �?                               @                              �?      @������R@33333�x@      �?              �?              F@      �?              �?                                       @       @      �?      �?        ������V@����L�@                      �?      �?     �P@      �?       @      �?       @       @       @               @       @       @                     P[@    ���@                                      8@      �?                                       @                                      �?      �?fffff�H@     E�@                                      �?      �?                                               @                              �?       @�����J@�����J@                      �?             @P@      �?               @      �?      �?      �?      �?      �?      �?       @                �����Y3@����̟�@      �?              �?      �?       @      �?              �?                       @               @       @              �?       @     �W@fffff��@                                      @      �?                                       @               @                               @fffff�L@fffff.d@      �?              �?             �Q@      �?       @      �?       @       @       @               @               @      �?       @     �X@�����R�@      �?              �?      �?     @Q@      �?       @      �?                       @               @       @              �?      �?������X@�����_�@                                      @      �?              �?                                       @                      �?       @      T@33333m@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?fffff&4@�����Q@      �?      �?                      .@      �?              �?                                               @              �?       @������S@fffff�@                                      ?@      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�4@     Z�@                                      �?      �?       @                                                                      �?        ������H@������H@                                     �N@      �?       @      �?       @       @       @       @       @       @      �?      �?       @fffff�]@3333�ż@      �?                              =@              �?                       @               @                                       @fffff&A@     f�@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @fffff�8@������@                      �?      �?      ?@      �?                       @               @       @       @       @      �?      �?      @�����IT@    ��@                                      >@      �?       @      �?               @                       @       @              �?       @�����Y@�����O�@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff�\@33333�@      �?                              8@      �?              �?                                       @       @              �?       @fffff�V@     }�@      �?              �?      �?     �P@      �?       @      �?       @                       @       @       @       @                fffff&Z@    ��@                                     �M@      �?       @               @       @       @       @               @      �?              �?fffff�S@������@                              �?     �D@      �?                                                                                        ������F@�����ǜ@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @                ����̜\@���̌��@                      �?      �?     �Q@      �?       @               @       @                       @               @      �?      �?�����LQ@����Y�@      �?                              9@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @     �4@fffff6@      �?              �?      �?      9@      �?              �?                               @       @                               @�����yU@����.�@      �?                      �?      D@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ffffff4@33333��@      �?              �?      �?      6@      �?              �?       @                                                                     �R@����̗�@      �?      �?                      �?      �?       @      �?                                                              �?       @����̬R@����̬R@      �?      �?      �?             @Q@      �?       @      �?               @       @                       @              �?        fffff�W@     �@              �?      �?             �P@      �?       @      �?               @       @               @       @      �?              �?fffff&Z@3333s��@      �?              �?             �K@      �?                       @       @       @                               @               @�����LM@33333��@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����9@�����F�@                                      1@      �?              �?                                                              �?       @     �Q@     �@              �?                      P@      �?       @                       @       @       @               @                      �?������R@����Y�@      �?      �?                      I@      �?       @               @       @                       @                      �?        fffff�Q@33333��@      �?                              E@      �?       @      �?               @                       @       @              �?       @     pY@3333s��@      �?                              "@      �?                                                                                      @�����yF@     �z@              �?                     �M@      �?       @      �?       @       @       @                                      �?       @     pV@ffff�x�@      �?              �?      �?      8@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @3333338@fffff�@      �?                              ,@      �?              �?                                       @       @              �?       @�����9W@������@      �?              �?      �?      F@      �?                               @       @       @                              �?      @33333�N@����ئ@      �?                              3@      �?                                               @       @                      �?      �?fffff�N@������@      �?              �?              P@      �?              �?       @       @               @       @       @       @      �?      �?33333Z@���̌͹@      �?                             �Q@      �?       @      �?       @       @       @       @       @       @      �?      �?        33333]@ffff�:�@                      �?             �J@      �?       @      �?               @                       @       @              �?      �?������X@    ��@                                      @      �?              �?                                       @                      �?      @33333T@�����u�@              �?                      �?      �?       @      �?                                                              �?      @����̜R@����̜R@                      �?              G@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?        33333s8@�������@                      �?              A@      �?       @      �?                                       @       @              �?       @�����iX@�����@                      �?      �?      R@      �?       @                               @               @       @       @      �?        333333S@3333s\�@                      �?      �?      I@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff&4@33333�@      �?              �?              G@      �?               @      �?      �?      �?      �?      �?      �?                       @������3@�������@      �?      �?      �?      �?      6@              �?               @                                       @                      @fffffD@�������@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @               @      �?      �?fffff�Z@�����|�@      �?                              "@      �?       @      �?                                       @                      �?       @fffffVU@����̴�@      �?                              E@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @����̌3@33333;�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?      �?              @33333�3@������G@      �?              �?      �?     �P@      �?       @      �?               @       @       @       @       @       @      �?        ������[@�����j�@      �?                              @              �?                               @                                      �?       @fffff�=@     �]@      �?                      �?      �?      �?                                                                              �?       @333333F@333333F@      �?      �?      �?              $@      �?              �?       @                                                               @33333�R@�������@      �?      �?                      @@      �?       @      �?                       @                                      �?      �?fffffFT@    �v�@                                      E@      �?                       @               @                                              �?fffffFK@����.�@      �?                      �?      6@      �?       @      �?               @                       @                      �?      �?fffffFV@�����u�@      �?                              2@      �?       @                               @       @       @       @      �?      �?      �?     �T@�����E�@      �?                              @      �?                                               @       @                      �?       @fffff�N@�����,o@      �?      �?      �?              �?      �?       @      �?                                                              �?       @������R@������R@                      �?      �?      D@      �?       @      �?               @       @               @                      �?      �?fffffX@����̖�@      �?                              :@      �?       @      �?                                               @              �?       @������T@fffff��@      �?                             �L@              �?               @               @               @       @              �?       @     �J@     ��@      �?      �?      �?              J@      �?       @      �?               @       @               @       @      �?      �?        fffffFZ@fffff �@      �?                      �?      @      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@fffff&M@                                     �F@      �?              �?       @       @                       @       @      �?      �?       @33333Y@3333�@                                      @      �?                       @       @                                                       @      L@�����Qx@      �?                             @P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?����̌3@�����
�@              �?                      @      �?              �?                                                              �?       @33333�Q@     pm@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @      �?        fffff&]@�����H�@                      �?             @P@      �?       @      �?               @       @       @       @       @       @      �?        ������Z@����٪�@              �?                      J@              �?                       @       @       @       @                      �?       @     @I@������@      �?                              ,@      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@     �q@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @     �4@33333Z@      �?                              @      �?              �?                                       @       @              �?       @�����V@fffff*w@      �?                              &@      �?                               @       @       @                              �?       @33333sN@     ��@                                     �@@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?33333�9@�����Љ@                      �?      �?      A@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        �����4@�����P�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@�����F@      �?                              P@      �?               @      �?      �?      �?      �?      �?      �?       @              @����̌3@�����`�@                      �?      �?     �Q@              �?               @       @               @       @       @       @              @33333SM@    @1�@      �?              �?              *@      �?       @               @                                       @              �?       @fffffvP@     2�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@������@@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����L4@�����L4@      �?                             �G@      �?               @      �?      �?      �?      �?      �?      �?       @                33333s4@     x�@      �?              �?             �G@      �?       @      �?               @       @       @       @       @              �?       @33333c[@���̌�@      �?              �?      �?     �Q@              �?               @               @       @       @       @       @                     �M@�����0�@                                      >@      �?       @               @               @               @       @      �?      �?      �?33333�S@33333��@      �?              �?      �?     �A@      �?       @      �?               @                       @                      �?        �����iV@33333��@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @33333�3@33333�3@                      �?      �?      3@      �?                                       @                                      �?        ������H@33333�@      �?      �?                      H@      �?       @      �?               @                       @       @      �?      �?       @     �X@����Y��@      �?              �?              E@      �?       @      �?               @       @               @                      �?             �W@3333��@                                      2@      �?       @               @               @                                      �?      @�����LN@fffff�@      �?                              @      �?                       @       @                                              �?        ������K@fffff�t@                                      5@      �?       @      �?               @                       @       @              �?      �?fffff�X@33333"�@      �?      �?      �?              =@      �?       @      �?                                               @              �?       @33333U@    �k�@      �?              �?              @      �?       @      �?               @               @                              �?       @�����YU@�����y@      �?      �?      �?      �?      I@      �?       @               @       @       @                       @       @      �?        ������R@ffff�ܭ@      �?                              3@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@fffffbv@      �?              �?      �?      @      �?                       @                                                      �?       @33333�H@fffffzr@                      �?              7@      �?       @      �?                       @                       @                      @������V@������@                      �?      �?      F@      �?               @      �?      �?      �?      �?      �?      �?                      @������3@     b�@      �?              �?      �?      .@      �?       @                               @       @                              �?        33333�M@������@      �?              �?             �N@      �?       @      �?               @       @               @       @              �?       @33333cZ@3333s��@      �?              �?      �?     �K@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �3@fffff	�@      �?              �?      �?      Q@      �?              �?       @       @               @               @       @                fffff�W@fffff�@                      �?             @P@      �?                       @               @       @                       @              �?33333sM@33333"�@      �?              �?              O@              �?                                       @       @               @      �?             �C@ffff�B�@                      �?      �?      7@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @������7@33333��@      �?                      �?      0@      �?       @               @       @                               @              �?       @fffffFQ@������@                      �?      �?      @      �?       @      �?               @       @               @                      �?      @33333�W@     6�@      �?              �?              =@      �?       @      �?               @                                              �?        �����	T@    ���@      �?              �?      �?     �I@      �?               @      �?      �?      �?      �?      �?      �?      �?              @ffffff3@     .�@                                     @P@              �?               @               @       @       @       @       @              �?������M@33333��@      �?                             @Q@      �?       @      �?               @               @       @       @      �?      �?        �����LZ@����ڼ@              �?      �?             �E@      �?       @      �?                       @       @       @       @      �?      �?       @33333�Z@ffff浱@                      �?      �?      ,@      �?       @      �?                               @       @                      �?       @������V@     T�@      �?              �?      �?     �M@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����L3@����̢�@                                      I@      �?              �?                       @       @               @       @      �?        �����lV@    �а@      �?              �?      �?      F@      �?       @       @      �?      �?      �?      �?      �?      �?      �?              @33333�9@     Z�@      �?                              .@      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@�����ys@      �?              �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              @33333s3@����̉�@                                      @              �?               @               @       @               @                      @      H@     Hi@      �?              �?      �?     �H@      �?       @      �?               @       @               @              �?      �?       @�����iW@ffff&��@      �?      �?                      "@      �?       @      �?               @                       @       @              �?      �?������X@33333��@                              �?       @      �?               @      �?      �?      �?      �?      �?      �?      �?                     �4@      C@                                      "@      �?              �?                                                                       @     �Q@fffff�@                      �?             �D@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�4@fffff\�@      �?                      �?      @      �?                       @               @                                              @33333�K@������c@                      �?      �?      3@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @������9@fffff^~@                                     �D@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������3@�����S�@                                      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @     @4@������Q@      �?              �?      �?      <@      �?              �?               @       @       @       @              �?                �����9W@3333���@      �?                              6@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     @9@     ��@      �?                      �?      �?      �?                                                                                       @      F@      F@                      �?      �?      1@      �?       @       @      �?      �?      �?      �?      �?      �?                      @�����8@fffff�y@              �?                      2@      �?       @      �?               @               @       @       @              �?      �?fffff�Y@fffff9�@      �?              �?      �?     �K@      �?                                       @       @                       @      �?      �?     �K@�����_�@                      �?      �?     �K@      �?                       @       @                                                       @������K@�����w�@      �?                              @      �?                                                                              �?        33333SF@     (t@      �?              �?      �?      @@      �?              �?                                                              �?             pQ@�����W�@              �?                      $@              �?                                       @                              �?       @fffff�=@fffff6r@              �?      �?              E@      �?       @      �?               @       @               @                      �?       @33333�W@33333��@      �?      �?                      @      �?               @      �?      �?      �?      �?      �?      �?                        �����4@������W@      �?                              J@              �?               @       @       @       @       @       @       @              �?33333�O@ffff��@      �?      �?      �?              @      �?       @               @       @               @                                       @�����P@     �}@                      �?              @@      �?               @      �?      �?      �?      �?      �?      �?                        ffffff3@33333	�@      �?              �?             �J@      �?       @      �?               @               @               @      �?                     pX@33333��@      �?              �?      �?     �J@      �?       @               @               @       @       @       @                       @�����lU@�����@                      �?              >@      �?       @      �?               @               @       @                      �?      �?fffff�W@ffff��@      �?                             �A@      �?               @      �?      �?      �?      �?      �?      �?                             �4@33333�@      �?                              @      �?                                               @                              �?      @ffffffI@�����Ii@                                      �?      �?              �?               @               @       @                               @������V@������V@      �?                              �?      �?       @                                                                              @     `I@     `I@      �?                              @      �?       @                                                                              @333333I@33333�i@                      �?      �?      8@      �?       @               @               @               @       @       @              �?fffff�S@�����ڜ@                      �?      �?     @P@      �?       @      �?       @       @               @       @               @      �?      �?33333�X@3333��@                                     �B@      �?       @      �?                               @       @       @                      �?33333Y@����̪�@      �?              �?      �?     �D@      �?                       @       @       @                              �?      �?        fffff&N@�������@                                     �A@              �?                                                                               @fffff&8@     d�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����4@�����4@                                      P@      �?       @      �?               @       @       @       @       @       @      �?      �?     �[@    @��@                      �?      �?     �F@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        fffff�8@33333ˑ@                                      @      �?              �?                                                              �?        33333cQ@������k@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @������3@������3@                                     �Q@      �?       @      �?       @       @       @       @       @       @       @              @33333�[@ffff�1�@      �?              �?      �?     �N@      �?              �?               @               @       @       @      �?      �?        ����̜X@33333�@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?ffffff4@fffff�Z@      �?                              M@      �?       @      �?                       @       @       @       @      �?      �?       @�����)Z@�����K�@                      �?      �?     �L@      �?                       @               @       @                      �?      �?      @fffff�M@3333���@                      �?               @      �?              �?       @                                                      �?       @������R@�����la@      �?              �?      �?      P@      �?              �?       @       @                                                       @33333CT@����Y�@      �?              �?      �?      L@      �?              �?               @       @       @                      �?      �?      @fffffvU@����̹�@      �?                               @      �?       @      �?                                                              �?       @fffff�R@������@      �?      �?              �?      L@      �?              �?       @                               @       @      �?              �?33333�W@����L��@      �?              �?      �?     �P@      �?       @                               @               @               @      �?        fffff�O@3333�]�@                                       @      �?              �?                                                                       @�����iQ@�����$b@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?       @33333�\@ffff�t�@      �?      �?      �?              @      �?              �?                                       @       @              �?       @     @V@������@      �?                              �?      �?              �?                                       @                      �?       @33333#T@33333#T@      �?      �?      �?              R@      �?                       @       @       @       @       @               @                ������R@    ��@      �?                               @              �?                                                                      �?      �?     @9@�����Ig@                      �?      �?      >@              �?                                       @       @       @                      �?������I@     f�@                                      �?      �?                                                                              �?       @33333�F@33333�F@                      �?              K@      �?       @      �?       @       @       @       @       @       @      �?      �?      @������\@    ���@                                     �C@              �?               @       @               @                      �?      �?        fffff&D@�����y�@                      �?      �?      1@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     �4@     $z@                              �?      ,@      �?                                       @               @                      �?      �?fffff�M@�����Ɖ@      �?              �?              A@      �?       @      �?                       @               @       @                       @fffff6Y@�������@                      �?      �?      @@      �?              �?               @                       @                      �?       @fffff�U@    �G�@      �?      �?                     �L@      �?       @      �?               @               @       @       @              �?        �����9Z@3333��@      �?              �?      �?      =@      �?                                       @       @       @       @       @              @33333�R@������@                      �?              J@      �?       @      �?               @       @               @                                fffff�W@����̡�@      �?                              8@      �?       @                                       @                      �?                �����LK@     i�@      �?                              �?      �?                       @                                                      �?      @�����YI@�����YI@      �?                              @      �?       @      �?                                               @              �?       @33333SU@����̌p@      �?              �?      �?      L@      �?                       @       @       @                               @      �?        fffff�M@ffff��@      �?              �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����Y4@fffffȖ@      �?              �?      �?      @@      �?              �?       @       @       @                       @      �?              @33333�W@����w�@      �?              �?              .@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������2@33333or@      �?              �?              D@      �?              �?               @       @                                      �?       @      T@    ���@                      �?              I@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ������3@�����x�@      �?                              F@      �?       @                       @       @       @       @       @      �?      �?             PU@����L�@                              �?      �?      �?       @       @      �?      �?      �?      �?      �?      �?                      @      8@      8@      �?              �?             �Q@      �?                       @                       @                       @                     @K@fffff��@      �?      �?                      R@      �?       @      �?       @       @       @       @       @       @       @                33333s\@����̥�@      �?                               @      �?                                               @                              �?      �?�����I@     P[@                                      N@      �?       @      �?               @       @               @       @       @               @�����,Z@����̽�@                      �?      �?      $@      �?       @               @       @                       @              �?               @33333�Q@33333!�@      �?                              @      �?       @       @      �?      �?      �?      �?      �?      �?                      @     @9@�����yY@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333s4@33333s4@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                      @�����Y4@     0W@      �?                      �?      @      �?                                               @                              �?        33333SH@ffffffm@              �?                       @      �?                                                                                       @������E@fffffFU@      �?              �?             �Q@      �?       @      �?               @       @       @       @       @       @      �?      �?fffff&[@ffff�
�@      �?              �?      �?      5@              �?                                                                      �?       @�����:@     ��@                      �?      �?      .@      �?               @      �?      �?      �?      �?      �?      �?      �?              @����̌4@33333r@                      �?      �?      @      �?                                               @                              �?      @ffffffH@������r@                      �?             �P@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?        ������4@�������@              �?                      �?      �?              �?                                                              �?       @ffffffQ@ffffffQ@                                       @      �?              �?                       @                                      �?       @33333�R@     d@      �?              �?      �?      ?@      �?                                       @       @                                      @�����,K@     ��@              �?      �?              L@      �?       @      �?                       @               @       @              �?        �����)Y@����8�@      �?              �?      �?     �I@      �?                       @       @               @                       @              �?     @N@ffff�b�@                      �?      �?      &@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @      9@33333�r@      �?              �?      �?     �N@      �?       @                               @       @       @       @       @      �?             @T@ffff&p�@      �?      �?                       @      �?               @      �?      �?      �?      �?      �?      �?                       @3333333@������B@      �?              �?              0@      �?              �?       @       @                                                             0T@33333��@      �?              �?      �?     �H@      �?                       @       @               @                                      �?������M@�����4�@      �?                              @      �?              �?               @                       @       @              �?       @     �W@     �@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              @������3@     "�@      �?                              (@      �?               @      �?      �?      �?      �?      �?      �?                      @33333s4@33333�o@                                      .@      �?       @               @                                                      �?      @������K@fffff�@      �?      �?      �?              @      �?              �?                                                              �?       @����̌Q@������q@                      �?              @      �?                                                                              �?      @�����G@�����D`@      �?                              �?      �?                                                                              �?      @������F@������F@      �?                              1@      �?       @      �?                       @       @               @              �?        ������W@     ��@              �?      �?              0@      �?       @      �?                                               @              �?      �?fffffVU@�����|�@      �?      �?                      �?      �?                                                                                       @������F@������F@                                       @              �?                                       @                              �?       @fffff�>@fffff�M@                      �?             @Q@      �?       @      �?       @                               @       @       @                ������X@����Yۺ@                      �?      �?     �I@      �?       @      �?                               @                              �?       @     0T@ffff��@                      �?      �?      R@      �?       @      �?               @       @       @       @       @       @      �?        �����L[@3333s�@                                      @      �?                       @                                                      �?       @������H@������s@      �?                              @      �?       @      �?               @       @               @       @                      @fffffZ@33333�@      �?                               @      �?              �?                                                              �?       @33333sQ@�����Tb@      �?              �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@fffff�3@                      �?      �?      @      �?       @                                                                      �?      �?�����yH@     q@                      �?             �N@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����L9@�����K�@                      �?      �?      9@      �?               @      �?      �?      �?      �?      �?      �?      �?              @�����4@�����@�@      �?              �?      �?      &@      �?               @      �?      �?      �?      �?      �?      �?              �?       @33333s4@�����Yo@                      �?      �?      7@              �?               @                       @                       @              @�����LA@�����k�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�3@fffff�3@                              �?      D@      �?                       @                       @       @                      �?      �?fffffP@3333�8�@              �?                      L@      �?       @      �?       @       @       @               @       @      �?               @     �[@    ���@      �?      �?                      �?      �?       @      �?                                                              �?       @     �R@     �R@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @3333334@������^@      �?              �?      �?     �J@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @ffffff3@fffffY�@      �?      �?                     �E@      �?       @      �?                                       @                      �?       @fffff6U@33333{�@      �?                             �O@      �?       @      �?               @                               @      �?              �?����̜V@    ���@      �?                              J@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@33333�@                      �?              M@      �?       @                       @               @                       @      �?      �?33333�M@33333b�@                      �?      �?      ?@      �?       @      �?                       @       @       @       @              �?       @�����Z@ffff�V�@              �?      �?              P@      �?              �?       @       @       @                       @      �?                     @X@ffff��@                      �?      �?       @      �?       @                       @                                                       @     �K@������{@      �?                              8@      �?                                               @                              �?      �?����̌I@fffff֓@      �?              �?      �?      Q@              �?               @       @                       @              �?              @ffffffF@����LO�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?                        fffff�4@33333cW@                                      @      �?       @      �?       @                                                      �?       @�����	T@������s@      �?              �?      �?      9@      �?               @      �?      �?      �?      �?      �?      �?      �?               @fffff�3@33333�@                                      I@      �?               @      �?      �?      �?      �?      �?      �?       @              �?ffffff3@�������@      �?                      �?     �C@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @      9@�����b�@      �?                              6@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����L4@fffff2}@                                      Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                     �9@33333w�@              �?                      "@      �?              �?                       @                                              �?     �R@33333�@              �?      �?      �?      @@      �?       @      �?                       @               @                      �?      @fffff�V@������@                                      �?      �?              �?                                                                      @fffff�Q@fffff�Q@              �?                      >@      �?       @      �?               @       @               @       @              �?       @fffffZ@33333b�@      �?              �?      �?     �G@      �?       @               @       @       @       @       @       @       @      �?      @     �V@����Yް@                                     �P@      �?       @               @       @       @       @       @       @       @      �?      �?33333�V@3333�M�@      �?      �?                     �C@      �?       @      �?                                       @       @              �?        ������W@����^�@      �?      �?      �?              R@      �?       @      �?       @       @       @       @       @       @              �?      �?�����9\@    �}�@                                      @      �?       @      �?               @       @       @       @       @              �?      �?�����y[@������@                                      �?      �?                                                                              �?      @fffff�F@fffff�F@      �?                              @      �?              �?                       @       @       @                      �?      @fffffV@�����`p@                      �?      �?      @      �?                       @       @                                                      �?33333�K@������v@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @fffff�3@fffff�3@      �?                              9@      �?              �?                                                                      @����̼Q@fffff��@      �?              �?      �?     �A@      �?               @      �?      �?      �?      �?      �?      �?       @                     �4@����̺�@      �?              �?      �?      <@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?�����L4@33333~@                      �?      �?      .@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @     @9@������x@      �?      �?      �?             @P@      �?       @      �?       @                               @       @      �?      �?       @     0Y@ffff��@                      �?      �?      Q@      �?       @      �?       @               @       @       @       @       @      �?        33333C[@���̌T�@              �?                      9@      �?       @      �?       @       @                       @       @              �?      @33333�Y@fffffȤ@      �?              �?      �?      R@      �?       @               @       @       @       @       @       @       @      �?        33333�U@ffff&?�@      �?                      �?      �?      �?                                               @               @              �?      @fffff�M@fffff�M@      �?      �?                      "@      �?                                               @                                      @������H@fffff�{@      �?                              @              �?               @       @                                              �?      @������A@fffff�Z@              �?                       @      �?              �?                                                              �?        ����̌Q@������\@      �?                             @Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�3@fffffݕ@                      �?      �?      @      �?              �?                                       @                      �?       @�����,T@fffff�m@              �?      �?      �?     �P@      �?       @      �?               @       @               @       @      �?      �?       @�����9Z@3333s�@      �?      �?      �?              M@              �?                       @       @                       @              �?       @fffff�F@fffff��@                                      @      �?                       @                       @                                       @�����K@     Ds@                                      (@      �?       @      �?       @                                                      �?       @����̼S@�������@                                      �?      �?              �?                       @               @       @                       @������W@������W@      �?              �?      �?     �K@      �?                       @       @               @                       @                fffff�L@�����̧@                      �?      �?     �F@      �?       @               @       @       @       @       @                              @33333ST@33333��@                      �?              5@      �?       @      �?       @               @               @       @              �?       @������Y@fffff��@      �?              �?             �Q@      �?       @               @       @       @       @       @              �?                ������S@ffff昵@      �?              �?              F@      �?       @      �?       @               @                                      �?      �?333333U@3333�T�@      �?              �?              6@      �?              �?                       @               @                      �?             �U@������@      �?              �?      �?     �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @                fffff�8@�����Q�@      �?                      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?      �?      �?      @fffff&4@33333Q�@                                      I@      �?               @      �?      �?      �?      �?      �?      �?      �?                     �3@fffff�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      �?����̌3@����̌3@              �?      �?              R@      �?       @               @       @       @               @       @       @      �?      �?fffffU@ffff��@                              �?      9@              �?               @                       @                       @                fffff�A@�����c�@      �?              �?             @Q@      �?                       @       @       @       @       @       @       @      �?      @�����,U@ffff���@      �?              �?             �N@      �?       @               @               @       @               @       @              �?fffff�R@����Ly�@      �?              �?             @P@      �?       @      �?       @               @               @       @              �?       @     Z@3333�@                      �?              N@      �?              �?       @                       @       @       @       @      �?       @�����LX@    ��@                      �?              R@      �?               @      �?      �?      �?      �?      �?      �?       @                ffffff3@�����a�@                                      Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �4@�����C�@      �?                               @      �?              �?               @                                                       @����̼R@     �b@                      �?      �?      (@              �?               @                       @                      �?              �?33333�@@     �{@      �?              �?      �?      K@      �?       @                               @                       @       @              �?����̬O@33333��@              �?                     �L@      �?                       @               @       @       @               @                fffffvQ@     F�@                                      G@      �?              �?                       @                                      �?      �?33333�R@�������@      �?      �?      �?              =@      �?       @                                                                      �?       @������I@     ��@      �?                              3@      �?                                                                              �?             �F@������@                      �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @                     �3@�����}�@      �?                      �?     �J@      �?              �?       @       @       @                       @      �?               @������W@ffff欳@      �?              �?              R@      �?                       @       @               @       @       @       @      �?        fffff�S@    @y�@      �?              �?      �?      (@      �?               @      �?      �?      �?      �?      �?      �?       @                �����5@�����`p@                                     �K@      �?                               @       @                       @       @      �?      @     0P@33333B�@                      �?      �?     �H@      �?                               @       @               @       @      �?              �?     �S@fffff�@                              �?      @      �?                       @                       @               @              �?              P@�����,f@                                      N@              �?                       @                       @       @              �?       @ffffffI@����̦�@                              �?      (@      �?                                                                              �?       @fffffFF@�����	~@      �?                              �?      �?                                                                              �?      @33333F@33333F@      �?              �?      �?      1@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @fffff&9@������y@                                       @              �?                                                       @              �?       @�����YA@      O@      �?              �?      �?      Q@      �?                                       @       @       @       @       @      �?        �����<R@    @Y�@                      �?             �@@      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@������@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @     @4@ffffffB@                                      �?      �?                                                                                      @     `F@     `F@      �?      �?                      @              �?                               @                       @              �?       @33333�D@fffff�`@                                      >@              �?                                       @               @      �?      �?      �?�����,D@33333��@                                      ;@      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff&3@�����U@      �?                      �?      J@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?������9@     ڔ@      �?                             @P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?        �����9@     ��@                              �?      @      �?                       @                       @                              �?      @����̌K@�����Tc@      �?                              A@      �?                       @               @                              �?              @�����yL@     ��@                      �?              P@      �?       @      �?       @               @               @               @      �?      �?fffff�W@3333�<�@      �?                      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@     �4@      �?              �?             �N@      �?       @               @               @                       @       @      �?      @�����yQ@3333���@      �?                              �?      �?       @                               @       @                                      @fffffO@fffffO@              �?                       @      �?              �?                                                              �?       @ffffffQ@�����t`@                                      :@      �?       @      �?                                                              �?        ����̼R@����̫�@                                       @      �?       @      �?                                       @       @                        ������W@�����P�@                                     �M@      �?       @       @      �?      �?      �?      �?      �?      �?       @               @33333s8@fffffT�@                      �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @              �?     `]@������@                                     �L@      �?                               @       @       @       @               @              @     pQ@�����l�@      �?                              :@      �?       @      �?                               @                              �?       @      T@�����Q�@                                       @      �?              �?                       @                       @              �?      @����̌U@fffffVf@                      �?      �?     �A@      �?              �?       @               @       @       @       @              �?       @������Z@ffff�X�@      �?              �?      �?     �J@      �?                               @               @       @                              �?     @P@�����G�@      �?      �?      �?              @      �?       @      �?       @       @                               @              �?      �?����̬W@������@              �?      �?              F@      �?              �?       @       @               @                              �?       @�����IU@     ��@      �?                             �@@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y4@     ��@                                      L@      �?       @      �?       @       @                       @       @              �?      �?fffff�Z@3333��@                      �?              H@      �?              �?               @       @               @       @      �?      �?       @33333CX@3333�T�@              �?      �?             �O@      �?       @      �?               @       @               @       @              �?       @     �Y@fffffO�@      �?              �?      �?      R@      �?       @      �?       @       @       @       @       @       @       @                33333�\@ffff9�@              �?                     �P@      �?       @      �?               @                                              �?      �?�����T@����Yh�@      �?      �?      �?      �?      G@      �?       @      �?       @       @       @               @                      �?       @�����,Y@33333��@      �?                              0@      �?                                               @                              �?      @������H@     ��@      �?              �?             �Q@      �?       @      �?       @       @       @               @       @      �?      �?       @ffffff[@ffff&��@      �?              �?              B@      �?       @      �?                                       @       @              �?       @������W@fffff$�@                      �?      �?      R@      �?       @               @       @       @       @       @               @                �����T@33333R�@      �?                              5@      �?               @      �?      �?      �?      �?      �?      �?                      �?     �4@�����-y@                                      @      �?               @      �?      �?      �?      �?      �?      �?                              4@333333a@              �?                      :@      �?       @      �?               @                       @                      �?       @�����IV@����Lˡ@                      �?      �?     �F@      �?                       @               @       @       @       @       @      �?      @     @T@33333��@      �?                      �?     �L@      �?       @               @       @       @       @       @       @       @              @33333cV@����Y��@      �?              �?      �?     �Q@      �?       @      �?               @       @               @       @       @      �?             �Z@3333�+�@                                      @      �?                       @               @                                              �?fffff�K@fffff�r@      �?                              G@              �?               @               @       @       @       @       @      �?             `N@����̚�@      �?                              .@      �?       @      �?                                                              �?      @      S@fffff��@                      �?      �?      P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      @�����8@�����\�@      �?              �?              .@      �?              �?                                                              �?        fffff&Q@fffffR�@      �?                              G@      �?       @      �?       @                               @                      �?      �?�����IV@���̌��@                                      @      �?                                                                              �?      �?fffffF@�����Di@      �?              �?      �?     �A@      �?       @                                       @       @       @      �?      �?        �����\R@33333ʤ@                                      �?      �?       @      �?                                       @                      �?       @fffff&U@fffff&U@                                      G@      �?       @      �?       @       @                                                      @     U@33333�@                      �?              (@      �?                       @                       @                                        �����K@     ��@      �?                              <@      �?       @      �?               @       @               @       @              �?       @�����lZ@     G�@                                      �?      �?                                                                              �?      @�����9F@�����9F@                      �?      �?      R@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�3@33333��@                      �?      �?      O@      �?              �?               @       @               @       @              �?       @�����	Y@����L��@      �?                              "@      �?       @      �?                                       @                      �?       @     `U@�������@              �?                      �?      �?              �?                                       @                               @����̜S@����̜S@                      �?      �?     �C@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      @3333338@����̔�@                                      ?@      �?                               @       @       @       @       @       @              @������S@fffff��@                      �?      �?      ,@      �?              �?                                                                       @����̌Q@     Z�@                                      D@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ������4@fffffډ@      �?                               @      �?              �?                       @                       @              �?       @fffffvU@������d@                                     @P@      �?                       @       @               @                       @      �?      @������M@�����7�@                                      A@      �?       @      �?       @       @       @               @       @              �?      @33333s[@    ��@                                      =@      �?       @               @       @               @                                      @������P@fffff$�@      �?              �?             �B@      �?       @      �?                       @       @       @               @              @33333�W@ffff�	�@                      �?      �?      D@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff&4@�����J�@      �?                             �B@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?fffff&4@     ��@      �?              �?             �N@              �?               @               @       @       @       @       @      �?      @33333O@3333���@      �?      �?              �?      C@      �?       @      �?       @                                                      �?      @�����T@����L��@      �?                              A@      �?       @      �?               @       @               @       @              �?       @fffff�Z@    ���@      �?                              *@      �?              �?                                               @              �?       @fffff6T@�������@                      �?      �?      M@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?      �?     �8@�����g�@                      �?             �Q@      �?       @                               @       @       @       @       @      �?        �����T@    @�@      �?                              @      �?              �?       @                                       @              �?      @33333�U@33333�n@              �?                       @      �?       @                       @                                              �?      �?fffffFL@     �]@      �?              �?      �?      K@      �?              �?               @               @                       @      �?        ������S@����
�@      �?                              $@      �?              �?       @       @       @               @       @              �?       @�����Z@������@              �?      �?              R@      �?       @      �?               @       @       @       @       @       @      �?      �?33333�[@    @ʾ@              �?                      �?      �?              �?                                                              �?       @�����iQ@�����iQ@      �?              �?      �?     �Q@      �?       @               @       @       @       @               @      �?                fffff�S@3333�E�@      �?      �?              �?      &@      �?                               @               @                              �?       @fffffFK@     ʂ@                                      �?      �?              �?                                       @                               @33333�S@33333�S@      �?              �?      �?      @      �?       @      �?                       @               @       @                       @�����IY@fffffx@                                      @      �?                               @                                                      �?�����YI@������b@                                      �?      �?                                                                              �?      �?fffffFF@fffffFF@      �?                      �?      @      �?                       @                                                               @����̬H@�����tk@                      �?             �A@      �?                       @                               @              �?      �?        33333O@ffff�N�@      �?                              �?      �?                                                                                      @fffff�F@fffff�F@                      �?              @      �?       @      �?                                                              �?      �?fffff�R@     �l@      �?      �?      �?              3@              �?                       @       @                                      �?      �?fffff&A@33333	�@      �?                             �@@      �?              �?               @       @                                      �?      �?     �S@�����!�@                              �?      @      �?                                               @                              �?      @     �I@������q@      �?              �?              2@      �?       @      �?                                                              �?       @�����IR@�����g�@      �?              �?             @P@      �?       @      �?               @                       @                      �?        fffff�V@�����4�@      �?              �?      �?      E@      �?       @      �?       @                               @       @      �?               @fffffFX@    �a�@      �?                             �E@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333s:@33333X�@                      �?      �?     �H@      �?       @      �?                                       @       @              �?        ������W@3333��@      �?      �?                      Q@      �?       @      �?               @       @                       @              �?       @������W@33333g�@              �?      �?              J@      �?       @      �?       @       @       @               @       @              �?       @fffffF[@3333��@              �?      �?              N@      �?       @      �?               @       @               @       @              �?       @�����yZ@    @�@      �?              �?      �?      R@      �?       @      �?       @               @               @       @       @      �?        33333cZ@    @v�@      �?              �?      �?      Q@      �?              �?       @               @                               @              �?fffffT@ffff&��@                      �?             �P@      �?       @      �?               @       @               @       @      �?      �?        �����lZ@3333�@                      �?             �H@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        fffff&4@�����j�@                              �?      1@      �?       @                               @                              �?      �?      @������K@     L�@      �?      �?                       @      �?                       @               @               @                                ������P@33333�W@      �?                             �F@      �?       @      �?       @               @       @       @       @              �?      �?�����[@3333�d�@              �?      �?             �B@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@fffff��@      �?      �?      �?             �Q@      �?       @      �?               @       @               @       @      �?      �?       @333333Z@3333�@      �?              �?      �?      ?@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @     �9@����̜�@      �?      �?                      @      �?       @      �?               @       @               @       @              �?       @     @Z@33333gr@                                      @      �?       @      �?                                                              �?       @     �R@33333�k@                                      &@      �?       @      �?       @                                                      �?             �S@fffff
�@                      �?      �?      2@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����9@33333�z@                      �?      �?      9@              �?               @       @       @               @       @              �?      �?�����LM@�����z�@                      �?              R@      �?       @      �?       @       @                               @       @      �?      �?����̜W@3333�	�@      �?                              ,@      �?              �?                       @                                               @�����S@33333v�@      �?              �?      �?      9@      �?       @       @      �?      �?      �?      �?      �?      �?              �?        ffffff9@������@              �?      �?              &@      �?              �?                               @       @                      �?       @������T@fffff��@      �?                              �?      �?       @               @       @                                                       @33333�N@33333�N@              �?      �?              Q@      �?       @      �?       @       @                               @      �?      �?      �?33333#X@ffff浹@                      �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�3@fffff��@      �?              �?             �J@      �?       @      �?       @               @                       @                       @�����yW@33333��@      �?              �?              ,@      �?       @      �?               @       @                                      �?       @������T@     ��@                      �?              @      �?               @      �?      �?      �?      �?      �?      �?                      @������4@      R@                      �?             �D@      �?              �?               @       @       @                      �?      �?        ����̌U@�����@      �?              �?             �M@      �?       @               @                       @               @      �?      �?      @fffffFQ@ffff� �@                      �?              R@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?      9@������@      �?                             �P@      �?       @       @      �?      �?      �?      �?      �?      �?      �?                33333s9@�������@              �?      �?              E@      �?              �?       @                                                      �?      �?������R@�����:�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @������3@������3@                      �?              0@              �?                                       @       @       @              �?       @������H@�����Q�@                      �?             �F@      �?              �?                               @       @       @       @      �?      �?������W@����̽�@                              �?     �H@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?33333s3@fffffʌ@                                     �D@      �?               @      �?      �?      �?      �?      �?      �?       @              @      4@fffffR�@                      �?             �Q@      �?       @               @       @       @       @       @       @       @              �?     pU@�����O�@      �?              �?              E@      �?       @               @                       @       @       @      �?              �?�����T@�����_�@              �?      �?              :@      �?       @      �?               @       @                       @              �?       @fffffvW@������@                                      R@      �?       @      �?       @       @       @       @       @       @       @      �?       @������\@����Y��@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?      �?               @����̌4@������X@                      �?      �?     �D@      �?       @      �?       @       @                       @                      �?        33333�W@33333k�@      �?      �?      �?              B@      �?       @      �?                                               @              �?      �?     PU@    �y�@      �?                              �?      �?              �?                                                              �?       @33333cQ@33333cQ@                                      *@      �?       @      �?       @                               @       @              �?       @fffffY@fffff;�@                                     �F@      �?       @      �?                       @       @                              �?       @     �U@fffffˮ@      �?                      �?      �?      �?              �?                                                              �?       @������Q@������Q@      �?                              6@      �?       @      �?               @                                              �?       @fffff�S@fffff	�@      �?                              @      �?                       @               @       @       @       @       @      �?      @     T@fffff�~@      �?                             �D@      �?              �?               @               @       @              �?      �?       @33333cV@    �#�@                      �?      �?      @      �?              �?               @               @                              �?       @      T@�����)n@                      �?             �Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?�����3@�����q�@                      �?      �?     �I@      �?       @      �?                       @                       @      �?      �?       @������V@�����ʱ@                                      �?      �?                                                                                      @����̬F@����̬F@                      �?      �?     �D@      �?                       @       @               @       @       @       @               @����̜S@ffff�l�@      �?                              G@              �?                       @                                                        �����L>@fffff��@              �?      �?              �?      �?              �?                                                              �?      @����̜Q@����̜Q@      �?      �?                     �A@      �?       @      �?       @                                       @                      �?     �V@     ٨@                      �?              9@      �?                       @       @               @               @              �?      @33333�Q@����̶�@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?              �?       @fffff�3@fffff�3@                      �?      �?      @      �?       @                       @       @               @                      �?        �����IQ@     `m@              �?      �?      �?     �N@      �?       @                               @               @              �?      �?       @�����LP@������@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      �?33333s4@fffff�T@      �?      �?      �?             �M@              �?               @               @       @       @       @       @      �?      �?33333P@3333�]�@      �?                               @      �?              �?                       @               @       @              �?       @fffff�W@fffff�h@                                      :@      �?              �?       @               @       @                      �?      �?      �?������U@33333ġ@      �?              �?              >@      �?       @      �?                                       @       @              �?      �?33333�W@ffff�d�@                      �?      �?      �?      �?              �?                                                              �?       @33333sQ@33333sQ@      �?                              @      �?              �?                                               @              �?       @������S@�����Dt@      �?              �?      �?      R@      �?       @               @       @       @                               @              �?�����P@     p�@      �?              �?              @      �?       @      �?                               @                              �?        ������S@     xo@                      �?              ,@      �?       @               @                               @                      �?        �����,P@     h�@      �?                      �?      5@      �?       @      �?       @                                                               @fffffT@�����L�@      �?              �?      �?      2@      �?                       @               @       @       @       @                       @     �T@�����,�@      �?              �?      �?     �N@      �?                       @       @       @       @       @       @      �?                �����9U@    ���@                      �?             �M@      �?       @      �?               @                       @       @                       @fffffFY@ffff旷@      �?              �?             �M@      �?       @      �?                       @               @       @      �?      �?             �X@����I�@                      �?      �?      =@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����:@fffff��@      �?                              ;@      �?                       @                                                              @�����,I@fffff�@      �?              �?              N@      �?       @      �?               @       @               @       @      �?                     �Y@������@      �?      �?                      4@      �?              �?                                       @       @                       @�����|V@�������@      �?              �?              F@              �?                       @       @               @       @       @                fffff&K@ffff欢@                                      C@      �?       @               @       @       @                                      �?        ������P@����̴�@      �?      �?                      &@      �?              �?                                               @              �?       @     �S@�����Q�@      �?              �?      �?      @      �?       @      �?       @               @                                      �?       @      U@     \|@      �?      �?                      "@      �?       @               @                                                               @fffffFK@������~@      �?      �?      �?      �?     @P@      �?       @      �?       @       @                                              �?       @     pU@3333s8�@                                      ?@      �?       @      �?                                                              �?       @33333S@�����g�@      �?                              @      �?              �?                                       @                      �?      @fffffT@������x@                              �?      �?      �?                       @                       @                                       @     @K@     @K@                                      @      �?       @                                       @       @                      �?       @������O@�����tc@                      �?              R@      �?       @      �?       @       @       @       @       @       @       @      �?             �\@    `<�@      �?                              :@      �?                                               @       @              �?              �?������M@     ��@      �?      �?      �?              D@      �?       @      �?       @                               @       @                       @fffffvY@������@      �?                              @      �?              �?       @                                                              @fffff�R@����̬�@      �?                      �?      1@      �?                                                                      �?              @�����LF@33333K�@                                      4@      �?       @                       @               @               @              �?      �?�����9Q@fffffi�@      �?              �?      �?      N@      �?       @      �?       @               @               @              �?      �?        ������W@     ��@                      �?      �?     �N@              �?                       @       @       @       @       @       @      �?        ������N@����LN�@      �?              �?              N@      �?                       @                               @              �?      �?      @fffff�M@����Lҫ@                                      ?@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�4@����̊�@                      �?              M@              �?               @       @                       @              �?      �?       @����̬F@33333أ@      �?                              �?      �?              �?                                       @                      �?       @     �S@     �S@      �?                      �?     �P@      �?                               @       @       @       @       @       @      �?      �?     �S@����L�@                      �?      �?      :@      �?               @      �?      �?      �?      �?      �?      �?       @              �?fffff�3@fffff�~@                      �?      �?      P@      �?       @      �?               @       @       @       @       @      �?      �?       @������[@3333�b�@      �?              �?             �O@      �?                       @       @               @       @              �?              �?33333�Q@�����`�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @     �3@     �3@                      �?      �?     @Q@      �?       @      �?               @       @       @       @       @      �?      �?             0[@����E�@      �?                              ?@      �?       @      �?               @                                              �?       @�����T@33333��@              �?                     �P@      �?       @      �?       @                               @       @       @      �?        ������Y@�����G�@              �?      �?              E@      �?       @      �?                                       @       @              �?       @33333�W@     Ѯ@                                      �?      �?                                                                                       @fffff�E@fffff�E@                      �?               @      �?               @      �?      �?      �?      �?      �?      �?                        fffff&4@     �c@      �?                              1@      �?       @      �?       @       @       @       @       @                      �?        ������Z@fffff �@      �?                             �J@      �?               @      �?      �?      �?      �?      �?      �?       @                fffff�3@     ��@      �?      �?      �?              @@      �?       @      �?                                               @              �?       @     @U@������@      �?                              M@      �?                               @       @       @       @               @                fffff�Q@ffff桯@      �?                              7@      �?       @      �?                       @                                      �?       @     @T@fffff��@      �?              �?              B@      �?              �?       @                               @       @              �?       @ffffffW@����L�@              �?                      7@      �?       @      �?                       @                                      �?      @fffff�S@33333��@      �?              �?      �?      =@      �?              �?                                                              �?       @     �Q@33333۞@      �?              �?      �?     �I@      �?       @      �?               @               @                      �?                �����U@    �˰@                      �?      �?      (@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?     @9@33333+q@                              �?      F@      �?       @                       @                       @       @      �?      �?      @33333cS@33333�@      �?                             �B@              �?                                               @               @              �?fffff�A@�������@                                       @      �?       @      �?               @                                                       @33333�S@     �b@                                      6@      �?                       @                                                      �?       @fffff�H@33333d�@                              �?      G@      �?       @      �?                       @       @                              �?        333333U@3333��@      �?                              7@      �?       @      �?                                                              �?       @����̼R@����̹�@      �?                              4@      �?       @               @                       @                                        ������M@����̜�@      �?                              Q@      �?              �?               @       @                              �?              �?fffff�S@3333sU�@                                      "@      �?                                                                              �?       @     �E@33333[y@                      �?      �?      ,@      �?              �?               @               @               @              �?      �?�����iV@fffff�@                      �?             �Q@      �?       @      �?                       @       @       @       @       @      �?        33333Z@    ��@      �?              �?      �?     �O@      �?               @      �?      �?      �?      �?      �?      �?       @              @����̌3@fffffv�@                      �?              .@      �?       @                                                                      �?       @����̌I@333339�@                                     �@@      �?              �?                                                              �?        ������Q@33333̢@      �?      �?      �?             �L@      �?       @                       @       @               @              �?      �?      �?fffff�Q@����,�@      �?                              E@      �?       @      �?                       @                                               @������S@������@                      �?      �?      @      �?                                                                                      @ffffffF@fffff�k@                                     �A@      �?       @      �?       @       @       @       @       @       @       @      �?      @�����L\@������@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                             �3@     �3@                      �?      �?      H@      �?       @      �?                                               @      �?      �?      @33333�T@ffff�{�@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �4@     �4@                                      @      �?                       @                       @                                      �?������J@�����<p@              �?      �?              N@      �?       @      �?                       @               @       @      �?      �?      �?      Y@     ��@                                      @@      �?       @      �?       @               @       @       @       @      �?      �?        33333c[@     0�@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �3@������q@      �?              �?      �?      =@      �?                       @                                       @              �?      @�����N@�������@      �?                              B@      �?       @      �?                                               @              �?       @�����9U@fffff��@      �?                              3@      �?       @      �?                                               @              �?             �U@������@                      �?      �?      8@      �?       @               @       @       @                               @               @fffffP@�����Z�@      �?                              C@      �?       @               @       @       @       @                                       @�����|Q@����ä@                      �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����9@fffff�@                      �?             �K@      �?       @      �?               @       @               @       @              �?      �?������Y@ffff�,�@                      �?             �A@      �?              �?                                                              �?       @33333�Q@�����@                      �?              D@      �?       @      �?       @               @               @       @      �?                     pZ@���̌��@      �?                              �?      �?              �?                                                              �?       @33333�Q@33333�Q@                      �?              H@              �?                       @       @                              �?              @�����YA@     �@      �?              �?              &@      �?                                                       @                      �?        fffff�K@33333�@      �?              �?      �?     �Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?        ������3@����̭�@                      �?      �?     �A@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @������3@������@              �?      �?              R@      �?       @      �?       @                                               @                     �S@    @�@                      �?             �D@      �?       @      �?       @       @       @       @       @       @              �?        ffffff\@3333��@      �?                             @Q@      �?       @               @       @       @       @       @       @       @              @������V@������@      �?                              @      �?                                                               @              �?      @fffff�K@     �m@                      �?      �?      ,@      �?       @      �?                       @                       @              �?       @     �U@fffff��@      �?              �?      �?     �B@      �?              �?                                       @       @      �?              �?������V@����_�@      �?      �?      �?             �Q@              �?               @       @       @       @                       @              �?�����,G@�����2�@      �?              �?      �?      *@      �?                               @       @       @                                        fffff�N@�����p�@                      �?             �I@      �?              �?       @       @       @               @              �?      �?       @     `W@���̌�@      �?                      �?      <@      �?              �?       @                                                      �?        ������R@����)�@      �?                      �?       @      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@33333sE@                                      �?      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @33333�9@33333�9@                      �?      �?      K@      �?                       @               @       @               @       @                �����|Q@3333�?�@      �?      �?      �?             �L@              �?                                               @       @              �?       @�����lF@ffff��@                      �?      �?      5@      �?                                                                              �?       @�����yF@     �@      �?              �?      �?     �B@              �?               @       @       @                                                �����D@33333��@      �?              �?      �?      <@              �?               @               @       @       @              �?              @ffffffI@33333��@      �?                              1@              �?                                                                      �?      @fffff�9@33333�{@                                      5@              �?               @                       @                       @              @����̌A@33333�@                      �?      �?      ,@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @33333�3@fffffzp@      �?                              3@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������2@33333sq@      �?                             @Q@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @�����3@fffffӓ@      �?              �?      �?      A@      �?       @      �?               @                       @       @              �?        �����lX@     ��@      �?              �?      �?      "@      �?              �?                       @       @       @       @                       @fffff�Y@�����S�@              �?      �?              :@      �?                                       @                       @      �?              @�����YN@�������@      �?                              $@      �?       @      �?       @                               @       @                       @33333�X@fffff��@              �?      �?              R@      �?       @               @       @       @       @       @       @       @      �?        fffffvV@����Y)�@              �?      �?             �P@      �?       @      �?       @               @               @       @      �?      �?      �?33333�Z@    ��@      �?      �?                      @              �?                       @               @               @              �?       @333333F@����̜p@                      �?      �?      R@              �?               @       @       @       @       @       @       @      �?      �?�����LP@3333s��@      �?                      �?      H@      �?       @               @       @       @                              �?      �?        �����P@3333���@                                     �G@      �?       @               @               @       @                       @      �?      @     @P@������@                                      �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff&3@fffff&3@                      �?      �?      6@      �?              �?                                               @              �?       @�����	T@�������@      �?                             �M@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����Y3@fffff.�@      �?                              "@      �?       @                                                       @                      @33333�M@33333�@      �?              �?             �O@      �?       @                               @       @       @       @       @              �?33333�S@������@                                       @      �?                               @                                              �?      @������H@����̬\@      �?                             �J@      �?                                       @                       @      �?      �?       @����̌N@�����;�@      �?                               @      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@������@@      �?              �?      �?     �A@      �?       @      �?               @       @       @       @       @              �?       @�����|[@����̌�@                      �?              R@      �?       @      �?       @       @       @               @       @       @      �?      �?������[@ffff���@              �?                      �?      �?              �?                       @                                      �?        33333�R@33333�R@                                      (@      �?              �?                       @       @               @              �?       @�����YV@������@      �?              �?      �?      M@      �?       @      �?               @               @       @              �?      �?      �?����̬W@����Y6�@                      �?      �?     �Q@      �?              �?                       @                               @               @33333S@3333s<�@      �?                              B@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?����̌2@     ��@                      �?              D@      �?               @      �?      �?      �?      �?      �?      �?       @              @�����3@�����`�@      �?      �?      �?             @P@      �?       @      �?               @       @               @       @              �?       @fffffZ@���̌��@      �?              �?      �?      N@      �?              �?               @       @               @              �?               @����̼V@fffffM�@                      �?              R@      �?       @      �?       @               @       @       @       @       @      �?      �?������[@33333ɾ@              �?      �?      �?      &@      �?       @      �?                       @                                      �?      �?fffff�S@������@      �?              �?              M@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@����̇�@                                      (@      �?       @                                       @       @       @      �?      �?      @fffff�R@�������@      �?                              @      �?                       @                       @                              �?      @     �K@33333�p@                                      R@      �?       @      �?                       @       @       @       @       @      �?      �?     �Z@3333���@                      �?      �?      4@      �?       @               @                               @       @      �?                      S@     Ә@              �?                     �Q@      �?       @                       @       @       @       @               @      �?             �R@ffff�\�@      �?                              $@      �?              �?                                                                      @������Q@     ��@      �?              �?             �H@      �?              �?               @                       @                      �?      �?33333SU@3333�ɰ@                                      H@      �?                       @       @                                       @              �?     �K@3333���@                      �?      �?      Q@      �?       @      �?               @               @       @       @       @      �?      �?     �Y@3333s�@                              �?      &@      �?               @      �?      �?      �?      �?      �?      �?                      �?33333�3@fffffk@      �?      �?      �?              G@      �?              �?                                               @              �?       @�����T@fffff*�@                      �?      �?     @P@      �?                       @       @       @                              �?                ����̬N@33333D�@                                      2@              �?                               @       @                              �?       @������A@fffff��@      �?                              6@      �?       @       @      �?      �?      �?      �?      �?      �?              �?      �?������8@fffff�~@                      �?      �?      ,@      �?                       @       @               @                                        ������M@�����f�@                      �?      �?      O@      �?       @      �?       @                               @       @       @      �?        �����IY@����Y�@                                     �K@      �?              �?               @       @                                      �?       @33333cT@    ���@                              �?     �P@      �?       @      �?       @               @       @                       @      �?      �?����̼V@����*�@      �?              �?              J@      �?       @                       @               @                                        ����̬N@����è@                      �?      �?     �O@      �?       @      �?       @                               @       @      �?      �?      �?������X@33333��@                                      @      �?               @      �?      �?      �?      �?      �?      �?      �?              @fffff�3@����̤e@                      �?              E@              �?                       @               @                      �?              @fffff�@@33333��@              �?      �?              @      �?       @      �?                                               @              �?       @33333#U@�����6�@                                      7@      �?              �?               @               @                              �?      @fffff�S@     ߛ@                      �?      �?      L@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      �?������3@������@      �?                              G@              �?               @               @       @                       @              @      C@fffffm�@      �?              �?      �?      0@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@�����(r@      �?                              $@      �?              �?       @       @       @       @       @       @              �?       @fffff�[@33333M�@      �?              �?      �?      P@      �?       @      �?       @       @       @                                      �?       @33333�V@    �H�@              �?      �?              <@      �?       @      �?               @       @       @       @       @              �?       @fffff�[@������@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                       @33333s3@33333s3@                      �?      �?     �E@      �?               @      �?      �?      �?      �?      �?      �?      �?              @      4@�������@                                      K@      �?       @      �?                               @       @       @              �?       @fffffY@ffff�@�@              �?                      4@      �?              �?                                       @                                �����,T@�����8�@      �?                              @      �?       @      �?               @                                                       @����̜S@����̠t@      �?              �?      �?     @P@      �?                       @                       @       @       @       @      �?        33333�R@ffff&Բ@              �?      �?      �?     �K@      �?       @               @               @       @       @              �?               @     S@���̌:�@      �?              �?      �?      J@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @����̌8@33333̔@                                      Q@      �?               @      �?      �?      �?      �?      �?      �?       @              �?������3@�������@              �?                      @      �?              �?               @       @               @       @              �?      �?33333�X@������{@                      �?      �?     �E@      �?       @      �?                       @               @       @              �?        33333�X@3333�q�@      �?      �?                      �?              �?                               @                       @              �?       @33333�C@33333�C@      �?                              $@              �?                                                       @              �?      @33333�@@33333�r@      �?                              @              �?                                       @               @              �?       @fffffD@fffffNd@                                      0@      �?       @      �?                                                                       @�����)R@33333��@                                      R@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     @4@�����{�@              �?      �?              K@      �?       @      �?       @       @       @       @       @       @      �?      �?        fffff�\@�����@      �?      �?                     @P@      �?              �?               @       @               @       @              �?        fffff�X@ffff&`�@                      �?      �?      I@      �?              �?                       @       @       @       @      �?              @33333�Y@    �!�@      �?              �?             @Q@              �?                       @       @       @       @       @      �?      �?      �?ffffffN@fffff��@              �?                      L@      �?       @      �?               @       @       @       @               @      �?        ������X@����LJ�@                                      �?              �?                                                                      �?      @fffff&9@fffff&9@      �?              �?      �?     �Q@      �?                       @       @       @               @       @       @      �?      �?�����	T@ffff&�@                      �?             �M@      �?       @      �?       @       @                       @                      �?       @     �W@ffff�ݵ@      �?              �?      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������4@     ��@                      �?             �B@      �?       @               @               @       @                      �?              �?fffffQ@    �^�@                      �?      �?      6@      �?                               @               @                                       @33333�K@33333ؒ@      �?                              �?      �?              �?                                               @                       @      T@      T@      �?      �?      �?              <@      �?       @      �?               @               @       @       @              �?       @33333sZ@     l�@      �?                              <@              �?                                       @                              �?      �?�����>@�����V�@      �?                              J@      �?                       @               @                              �?               @     �J@����Lͥ@                                      ,@      �?              �?               @               @                              �?      �?33333T@33333a�@      �?      �?      �?              0@      �?       @      �?                                       @                      �?      �?33333CU@�������@                      �?      �?     �C@      �?                       @                                                              �?fffff�I@     $�@                      �?      �?      &@      �?                       @                                                                     �I@�����-�@                      �?      �?     �A@      �?       @       @      �?      �?      �?      �?      �?      �?              �?       @     �9@fffff��@      �?              �?      �?      M@              �?               @       @       @               @              �?              @      I@3333�Ϧ@                                      A@      �?                       @       @                               @      �?               @fffffP@����
�@      �?              �?              ?@      �?       @                                               @                      �?      �?fffff�M@33333k�@                                      (@      �?       @      �?               @                               @              �?       @�����IV@33333��@                                     �@@      �?       @      �?               @       @               @       @                       @33333�Z@     {�@      �?                              *@      �?              �?                                       @       @              �?       @fffff�V@����̾�@                      �?      �?      7@      �?              �?               @       @       @                                       @33333�T@     ��@      �?                      �?      �?      �?       @      �?                                                              �?       @fffff�R@fffff�R@      �?                              �?              �?                                                       @              �?             �A@     �A@              �?                     �Q@      �?       @      �?                       @               @       @       @                33333Z@���̌��@                      �?              7@      �?       @                                       @       @       @              �?      �?�����iR@     ��@      �?      �?      �?             �H@      �?                               @                                       @              @fffff�H@����̼�@      �?              �?      �?      C@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?�����9@������@                                      �?      �?               @      �?      �?      �?      �?      �?      �?              �?      @�����3@�����3@                                     �@@      �?       @               @       @                                              �?      @33333sN@fffffǟ@                      �?             �P@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?     @9@������@      �?              �?             @Q@              �?               @               @       @       @       @       @                      N@     ��@      �?              �?              @      �?               @      �?      �?      �?      �?      �?      �?              �?      �?����̌4@33333�I@                                      3@      �?       @                               @                                      �?      @�����L@�����'�@                                      @      �?       @      �?                                                              �?       @fffffvR@     �@      �?                              �?      �?              �?                                       @       @              �?       @�����yV@�����yV@                                      ,@      �?              �?               @                               @              �?       @33333�U@�����s�@                                      �?      �?              �?                                                                       @fffff�Q@fffff�Q@                      �?      �?     �C@      �?       @      �?                               @       @       @              �?      �?������X@�����n�@                                      *@              �?                                                                      �?       @fffff�7@������r@      �?                              �?      �?              �?                                                              �?       @fffff�Q@fffff�Q@                                      G@      �?       @      �?                                       @       @                        33333X@    �/�@      �?              �?      �?      F@      �?                               @               @                              �?        33333sK@33333�@                                      (@      �?       @                                       @       @       @      �?              @33333�R@33333E�@      �?                             �E@      �?       @      �?                               @       @       @      �?      �?       @      Y@���̌s�@                                      B@      �?       @      �?               @       @               @       @      �?      �?        333333Z@ffff�\�@      �?              �?      �?     �N@      �?              �?               @       @       @       @       @      �?              �?������Y@ffff&1�@                      �?      �?     �H@      �?       @                       @               @       @       @       @                33333�S@ffff�|�@                                     �M@      �?       @               @                       @               @      �?                �����,Q@ffff�ͯ@                                      @              �?               @       @               @               @                      �?�����yI@�����9s@      �?                             �M@      �?                                       @       @       @                      �?       @�����)P@ffff�.�@                                     �D@      �?       @      �?       @                                                      �?      �?33333ST@����L�@      �?                              @      �?       @      �?                                       @       @              �?       @fffff�W@fffff�@      �?              �?             �N@      �?              �?               @       @       @               @                      �?������W@�����c�@      �?              �?              R@      �?       @               @               @       @       @       @       @              �?������U@    @η@      �?                              ?@              �?                               @               @       @      �?      �?       @fffffI@�����͗@      �?              �?             �H@      �?       @      �?               @                       @       @              �?        33333�X@    ���@      �?              �?      �?     �J@      �?              �?               @               @       @                      �?       @33333#W@3333s��@              �?      �?             �I@      �?       @      �?       @                                                      �?       @     `S@3333���@      �?              �?      �?     �G@      �?              �?       @               @                       @                       @33333�V@33333)�@                      �?              G@              �?               @       @                       @                               @fffff�F@����L�@                      �?               @      �?                       @                                       @              �?      @33333O@fffffF\@              �?      �?             �J@      �?       @      �?                                       @       @      �?      �?      �?fffff�W@    @��@      �?                              @      �?       @      �?                       @               @                      �?       @����̜V@�������@      �?              �?              @@      �?       @      �?                               @                      �?      �?       @     �S@����Lv�@                              �?      H@              �?                       @       @                       @                      �?fffff�F@3333�x�@      �?              �?      �?     �L@      �?               @      �?      �?      �?      �?      �?      �?       @              @     �4@�������@                                      �?      �?              �?                                                                      @fffff�Q@fffff�Q@      �?                              9@      �?                       @       @               @       @       @              �?      @     �S@     ��@              �?                       @      �?              �?                                                                       @     �Q@33333[c@      �?                              @      �?                               @                                                      @     �H@fffffj@                      �?      �?     �K@      �?               @      �?      �?      �?      �?      �?      �?       @              @      5@33333�@      �?      �?      �?              B@      �?                                       @       @                      �?              �?�����K@fffff#�@                                      H@      �?              �?               @                                      �?               @������R@����Ly�@                                      K@      �?       @      �?               @       @       @       @       @                       @fffff�[@�����~�@      �?              �?             @Q@      �?       @      �?                       @               @       @      �?                     �X@3333s��@      �?              �?      �?     �O@      �?       @       @      �?      �?      �?      �?      �?      �?       @              �?fffff�8@     ��@      �?                             �Q@      �?       @               @       @       @       @               @       @                fffff&T@33333L�@                      �?              @              �?               @                                                      �?       @�����=@333333`@                              �?      G@      �?              �?       @       @               @       @       @      �?      �?        �����LZ@�����ֲ@                                      3@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?     @4@fffff�w@                      �?             �E@      �?       @      �?               @                                                       @�����T@����̍�@      �?                              �?      �?              �?                                               @                       @fffff�S@fffff�S@                                      @              �?                               @                       @                       @     �C@     Xj@      �?      �?                      *@      �?       @      �?               @       @               @       @              �?       @������Z@33333Q�@                      �?             �H@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?33333�4@33333 �@                      �?      �?      Q@      �?       @      �?                                       @              �?      �?       @     �T@�����5�@                                       @      �?              �?               @                                                       @fffff�R@fffff��@      �?              �?              J@      �?                       @       @                       @       @      �?      �?      @������R@ffff�2�@                      �?      �?      R@      �?       @               @               @       @       @       @       @              �?�����,U@ffff��@              �?                      ?@      �?              �?       @                                                      �?      �?33333cR@����L]�@                      �?      �?     �M@      �?       @      �?               @       @               @       @      �?      �?       @������Z@33333p�@      �?                             �I@      �?       @      �?       @       @                       @              �?      �?       @33333�W@������@              �?                      :@      �?       @                                       @               @              �?       @33333�P@�����љ@      �?      �?      �?      �?      C@      �?       @      �?               @                       @       @                       @�����IY@3333�;�@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @     �3@     �3@      �?              �?      �?      R@      �?       @      �?       @       @               @               @       @      �?      �?     pX@�����O�@      �?              �?      �?      M@      �?       @      �?                       @       @       @       @      �?      �?        33333CZ@�����t�@                                      .@      �?                               @                                                       @�����lH@fffff�@                                     �E@      �?       @                       @       @       @       @       @      �?              �?fffffFU@    ���@                                      *@      �?                       @       @               @               @                        33333�P@     R�@      �?              �?      �?     �Q@      �?              �?       @       @       @       @       @       @       @              �?33333S[@�����f�@      �?      �?                       @              �?                                                                      �?      @33333s8@     �G@                                      G@      �?                                                               @      �?              �?33333�K@3333��@                      �?             �P@      �?       @               @       @       @                       @      �?              @fffff�R@3333sȳ@      �?                             �H@      �?       @      �?                                                              �?        fffff�R@3333��@      �?              �?      �?      @      �?               @      �?      �?      �?      �?      �?      �?              �?             @4@fffff�e@      �?              �?      �?     �@@      �?               @      �?      �?      �?      �?      �?      �?      �?              �?�����4@fffffd�@                      �?      �?     @P@      �?       @               @       @               @       @       @       @      �?             �T@����_�@                                      @      �?              �?                       @                                      �?      @     �R@33333�m@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @ffffff4@ffffff4@                              �?      (@      �?       @      �?       @                                                      �?       @33333�S@     j�@      �?                              7@      �?              �?       @               @               @       @      �?      �?      �?������X@    ��@      �?                              7@      �?               @      �?      �?      �?      �?      �?      �?                       @������4@fffff�}@      �?              �?      �?      L@      �?       @               @       @               @               @       @      �?      �?fffff�R@33333��@      �?              �?      �?      Q@      �?              �?       @       @       @               @       @       @      �?      �?     �Y@fffff��@                      �?             �O@      �?       @      �?               @       @               @       @      �?      �?       @     �Z@    �ٺ@      �?                              �?      �?              �?               @                               @              �?       @     @U@     @U@      �?              �?      �?     �H@      �?       @      �?                                       @                               @      U@����ٞ�@      �?              �?              ;@      �?                               @               @                              �?       @fffff�J@fffff��@                      �?             �K@      �?       @      �?       @                               @                      �?        33333sV@�����_�@                                      D@              �?               @                       @       @       @      �?      �?        fffffFK@fffffx�@      �?                      �?      (@      �?       @      �?                                                              �?      �?     pR@33333;�@      �?              �?      �?     �Q@      �?                               @               @       @       @       @      �?      �?fffffVR@    �"�@      �?                              @      �?       @      �?                                       @       @              �?       @fffffvW@�����܃@                      �?      �?     �J@      �?               @      �?      �?      �?      �?      �?      �?      �?                ����̌3@33333�@                                     �B@      �?       @               @       @       @       @       @                      �?      �?������S@ffff�A�@      �?              �?              �?      �?              �?                                       @                      �?       @33333#T@33333#T@      �?      �?      �?             �C@      �?       @      �?               @       @               @       @              �?       @�����iZ@����̼�@                      �?      �?     �O@      �?               @      �?      �?      �?      �?      �?      �?       @              �?      4@     �@                                      J@              �?               @       @               @                       @              @����̌C@fffff��@              �?                      @@      �?                               @               @                                        33333SK@fffff��@      �?                              �?      �?              �?                               @                              �?      @33333�R@33333�R@      �?                              �?      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�2@fffff�2@      �?                      �?      1@      �?                       @                                                      �?      @fffff&I@fffffv�@                      �?      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333s9@fffffU�@      �?                             �Q@      �?       @      �?       @                       @       @       @       @      �?      �?      Z@ffff&R�@      �?                              R@              �?               @       @       @       @       @       @       @      �?        ������O@�����p�@              �?                      �?      �?              �?                                                              �?       @����̌Q@����̌Q@                      �?             �M@      �?              �?               @               @       @       @       @      �?      @33333Y@����ْ�@                      �?      �?     @Q@      �?               @      �?      �?      �?      �?      �?      �?       @              @ffffff3@������@                                      O@      �?       @      �?                                       @       @      �?      �?             �W@33333}�@                      �?             �P@      �?               @      �?      �?      �?      �?      �?      �?       @              @fffff�3@�����ܔ@                                      J@      �?                       @               @       @                      �?              �?������L@    �ħ@                      �?      �?     �Q@      �?       @      �?       @       @       @       @       @       @       @      �?      �?33333C\@������@                                      ,@      �?                                               @               @      �?              �?����̌M@�����&�@                      �?      �?      B@      �?       @               @       @       @       @       @       @       @      �?      �?�����9W@    �f�@      �?              �?      �?      @              �?               @                               @                              �?fffffFC@33333�c@      �?                              1@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333s3@�����w@                                     �K@      �?                                                                      �?                fffff�F@33333=�@      �?                      �?      @      �?       @      �?                               @                                      �?333333T@33333�t@              �?      �?             �P@      �?       @                       @       @               @       @       @      �?        33333#T@������@      �?              �?      �?      H@      �?       @      �?       @       @       @       @       @       @       @              �?33333�[@ffff�C�@      �?              �?              R@      �?                       @       @       @       @       @       @       @              @�����U@������@      �?                      �?       @      �?       @               @       @                                                        �����yN@33333�`@      �?                              8@      �?              �?                               @       @       @              �?       @      X@ffff攠@      �?              �?              K@      �?                       @       @                       @       @       @      �?        33333�R@3333s_�@      �?              �?      �?      R@              �?               @       @       @       @       @       @       @      �?      �?fffffFP@����L��@      �?              �?              0@      �?       @      �?                                                              �?       @������R@�������@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @      �?      �?        33333s]@fffff��@                      �?             �I@      �?       @      �?                       @               @       @      �?      �?       @fffff�X@���̌S�@                                      3@      �?                               @                       @              �?               @�����M@     U�@                                      B@      �?       @               @                                              �?              @�����9K@     ��@                                      9@      �?       @      �?               @                       @       @              �?       @     Y@    ���@                      �?             �Q@              �?                       @       @       @       @       @       @                fffff�L@�������@                                       @      �?                                                                              �?      @     �F@����̌R@      �?                              @@      �?               @      �?      �?      �?      �?      �?      �?      �?              @������3@�������@                      �?      �?      "@      �?               @      �?      �?      �?      �?      �?      �?      �?              @     @4@33333�e@                                      2@      �?       @      �?                               @       @       @              �?        fffff�X@�����Û@      �?              �?             �I@      �?       @      �?       @       @                               @      �?      �?      �?�����X@����/�@      �?                             �E@              �?                               @       @               @      �?               @33333F@33333-�@      �?      �?      �?              0@      �?              �?                       @       @               @              �?       @33333�V@33333�@      �?              �?      �?     �Q@      �?       @               @       @       @       @       @       @       @               @fffff�V@    @��@      �?                              @      �?                                               @                              �?      @      I@�����	c@      �?                              5@      �?               @      �?      �?      �?      �?      �?      �?                      @      4@33333z@                      �?      �?     �H@      �?                       @               @       @                                             �N@����L��@      �?                              G@      �?       @      �?               @       @               @              �?      �?      �?������W@3333�F�@      �?                      �?     �J@      �?               @      �?      �?      �?      �?      �?      �?       @                     �3@fffffq�@                      �?      �?     �G@      �?                               @               @               @       @                fffff�O@    �~�@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�4@     `[@      �?                              �?      �?                                                                              �?       @33333sE@33333sE@      �?                              G@      �?       @      �?                                                                        333333R@�����b�@      �?              �?      �?      ?@      �?       @      �?       @               @               @              �?                33333�X@33333�@      �?                              �?              �?                                                                      �?       @fffff&9@fffff&9@      �?      �?                     �A@      �?       @      �?                                       @       @              �?       @������W@����$�@      �?                      �?     �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @�����Y8@fffffڙ@      �?                              @              �?                       @                       @       @              �?      @     �I@33333s@                                      @      �?               @      �?      �?      �?      �?      �?      �?                       @     �3@�����lM@      �?              �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                33333s8@�����
�@                              �?      $@      �?       @               @               @       @               @      �?              �?33333cR@fffff��@      �?                      �?      �?      �?       @                                                                      �?       @fffffI@fffffI@      �?              �?      �?      @      �?              �?                                                              �?      @33333cQ@fffff�q@      �?                              @      �?       @                                                                                333333I@     (a@              �?      �?              I@      �?       @      �?                               @       @       @      �?      �?       @�����)Y@    �E�@      �?              �?             �G@      �?               @      �?      �?      �?      �?      �?      �?      �?                fffff�3@�����w�@                      �?             @Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?33333�8@fffffٚ@              �?      �?      �?      (@              �?                                       @                              �?      @�����L=@fffff>v@                                      @      �?               @      �?      �?      �?      �?      �?      �?              �?      @      4@������N@      �?                              M@      �?       @       @      �?      �?      �?      �?      �?      �?       @      �?      �?33333s8@fffff��@                                     �G@      �?              �?       @                                                              �?������R@33333��@                      �?              5@      �?              �?                               @       @                      �?       @33333�U@�����k�@      �?              �?              2@      �?                                                                              �?        �����,F@fffff �@                      �?      �?      7@      �?               @      �?      �?      �?      �?      �?      �?       @      �?      @fffff�3@�����8|@      �?                      �?     �@@      �?       @      �?       @               @                       @              �?        33333�W@����L��@      �?                              ;@      �?               @      �?      �?      �?      �?      �?      �?      �?                �����4@����̔�@                                      8@      �?       @      �?                       @               @                      �?      �?�����<V@    �1�@                                      @      �?                               @               @       @       @              �?       @33333�R@33333�n@      �?                              �?      �?                                               @                                      @fffff�H@fffff�H@              �?                     �E@              �?               @       @                                              �?      �?������@@     q�@                      �?      �?     �P@      �?               @      �?      �?      �?      �?      �?      �?       @      �?             @3@�����s�@                      �?              @      �?              �?                                       @                      �?       @fffffFT@33333�@                                      6@      �?                               @       @               @              �?                     PP@33333��@      �?                              �?      �?                                                                              �?      @������F@������F@                      �?      �?     �B@      �?       @      �?               @                       @                      �?       @333333V@�����@      �?                              5@      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�3@fffffz@                      �?             �Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @              @������7@fffff �@                                      1@      �?               @      �?      �?      �?      �?      �?      �?                      �?33333�3@�����Eu@                                     �P@              �?               @       @       @       @                       @      �?      @33333�G@    �Ҩ@                              �?      2@      �?               @      �?      �?      �?      �?      �?      �?      �?                fffff&4@�����mx@                      �?      �?      �?      �?               @      �?      �?      �?      �?      �?      �?                      @�����4@�����4@                                      @      �?                       @                       @       @                      �?       @fffffP@fffff
v@      �?              �?             �A@      �?       @      �?                               @               @              �?        fffffvV@fffff��@                                      @      �?              �?       @                                                      �?       @33333�R@�����4m@              �?                      @      �?       @      �?                       @                       @              �?       @fffff6V@33333Gw@      �?              �?      �?      R@      �?       @       @      �?      �?      �?      �?      �?      �?       @                �����L8@     ��@      �?                              K@      �?       @               @               @       @       @       @       @                fffff�U@33333�@              �?                      ,@      �?              �?       @       @                                                       @fffff�S@33333O�@                      �?             �Q@              �?               @               @       @               @       @      �?        ������H@fffffT�@      �?                              8@      �?                       @                                                      �?        fffff�H@������@                      �?      �?      7@      �?       @      �?                                               @                       @ffffffU@�����1�@      �?      �?                      @      �?              �?                                                                       @fffffVQ@fffffZp@      �?              �?              @              �?                                                       @              �?       @33333�A@     �X@                      �?              A@      �?                                               @                                        �����I@33333]�@                      �?      �?      N@      �?                               @       @       @       @       @       @      �?        fffff&T@3333�R�@      �?                              �?      �?              �?               @                                              �?       @fffff�R@fffff�R@                                      @      �?              �?               @                       @       @              �?       @fffff�W@fffff6s@      �?              �?      �?      @              �?               @       @       @               @       @                      @�����lM@33333}@                      �?              2@      �?                                               @                              �?      @fffff&I@     f�@              �?                      2@      �?       @      �?               @               @                              �?       @�����\U@fffff��@                                      9@              �?                               @       @       @       @      �?               @�����K@�����<�@      �?              �?      �?      R@      �?       @      �?       @       @       @       @               @       @      �?      �?�����9Z@ffff�4�@      �?                              @      �?                       @               @                                               @     `L@����̤n@      �?                             �I@      �?               @      �?      �?      �?      �?      �?      �?      �?               @�����3@fffff~�@      �?              �?             @P@      �?       @      �?       @       @       @                              �?               @     pV@�������@                                      �?      �?       @      �?               @                       @       @              �?      �?     Y@     Y@      �?                             �P@      �?       @      �?               @               @       @       @      �?      �?       @     Z@�����̺@                      �?      �?     �I@              �?                               @       @       @       @      �?      �?       @33333L@ffff楦@                      �?      �?      G@      �?               @      �?      �?      �?      �?      �?      �?       @              �?ffffff3@33333�@                                     @Q@      �?       @               @               @       @       @       @       @      �?      �?fffffVU@fffff	�@                                      1@      �?              �?               @                       @                      �?       @33333�T@�����Ĕ@      �?                             �K@      �?              �?       @       @                       @       @      �?      �?      @�����9Y@������@                                      @      �?               @      �?      �?      �?      �?      �?      �?                      @fffff&4@�����|]@                      �?      �?      A@      �?               @      �?      �?      �?      �?      �?      �?                      @fffff�4@33333c�@      �?              �?             �A@      �?                       @       @       @                                              @     �N@ffff椠@                                      8@      �?       @      �?                               @               @              �?       @33333cV@3333���@      �?              �?      �?      8@      �?                       @       @               @               @              �?      �?33333�Q@����̩�@      �?              �?      �?      3@      �?               @      �?      �?      �?      �?      �?      �?       @              @3333334@fffff6x@              �?                      @      �?              �?       @       @                                                       @�����,T@�����lw@                                       @      �?               @      �?      �?      �?      �?      �?      �?              �?        33333�4@������C@                      �?      �?      I@      �?       @                       @       @       @       @       @      �?      �?      �?�����	U@fffffD�@      �?              �?      �?       @      �?                       @                                                      �?      �?fffff�I@������y@      �?              �?      �?      Q@      �?       @       @      �?      �?      �?      �?      �?      �?       @                ffffff9@�����P�@      �?                              @      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�2@�����Q`@                      �?      �?     �P@      �?                                               @                      �?      �?      �?33333�H@3333�g�@      �?                              A@      �?                               @                                              �?       @fffff�H@������@                                      3@      �?       @      �?       @       @                               @              �?       @������W@     ��@      �?                              �?      �?                                                                              �?        ������E@������E@      �?              �?              R@      �?       @      �?       @       @       @       @       @       @       @              �?����̜\@ffff�[�@                      �?      �?      R@      �?                       @       @       @                       @       @              �?     0Q@33333�@      �?              �?      �?     �Q@      �?       @                       @       @       @       @       @       @      �?      �?�����|U@    �+�@                                       @      �?              �?                                                                       @fffff�Q@     ha@      �?              �?             �Q@      �?       @               @               @       @               @       @              �?33333SS@33333z�@      �?                              "@      �?       @      �?                                                              �?       @     S@�����f�@                                      B@      �?               @      �?      �?      �?      �?      �?      �?      �?              @����̌3@     f�@      �?                              1@      �?                       @       @                                      �?              @�����L@�������@                      �?      �?      P@      �?       @      �?       @       @       @       @       @       @      �?               @fffffV\@    �6�@      �?                             �J@      �?               @      �?      �?      �?      �?      �?      �?       @              �?     �3@     j�@              �?      �?              �?      �?                                                                                       @      G@      G@      �?      �?      �?              @      �?       @      �?                                       @       @              �?        fffff�W@�����"�@      �?                              Q@      �?       @      �?       @       @       @       @       @       @      �?      �?      �?�����L]@3333�c�@      �?                      �?      ;@      �?               @      �?      �?      �?      �?      �?      �?       @              �?33333�3@������@      �?      �?      �?              @      �?              �?               @                               @              �?       @�����U@333339�@                      �?             @P@      �?                       @               @                                      �?      @33333�K@����L��@              �?      �?              ?@              �?               @       @       @                       @      �?      �?      �?333333I@fffff��@                                      �?      �?              �?                                       @                      �?       @     T@     T@                      �?      �?      K@      �?       @       @      �?      �?      �?      �?      �?      �?      �?      �?             �8@�������@                      �?              @      �?              �?                                                              �?       @�����<Q@     �u@                      �?              @      �?       @      �?               @                       @                      �?       @������V@fffff�v@      �?              �?             �Q@      �?       @               @                       @       @       @       @      �?      �?�����<S@����̩�@      �?                             �D@      �?              �?                               @                              �?       @     �R@33333"�@              �?                      2@      �?               @      �?      �?      �?      �?      �?      �?      �?                �����Y4@�����w@      �?                              0@      �?               @      �?      �?      �?      �?      �?      �?              �?      @33333�3@ffffffu@                      �?              R@              �?               @       @       @       @       @       @       @                     `P@3333�7�@                      �?      �?     �N@      �?       @      �?       @       @       @       @       @       @       @              �?fffff�\@ffff&`�@�?       �t�b�n_samples_fit_�M:�_tree�N�_sklearn_version��1.2.2�ub.